module dds#(
parameter phase = 0
)(
input clk,
input [13:0]freq,
output reg signed [13:0]dds_o 
);


reg signed [13:0] sin_rom [0:1953];
initial begin
sin_rom[0] = 0;
sin_rom[1] = 26;
sin_rom[2] = 52;
sin_rom[3] = 78;
sin_rom[4] = 105;
sin_rom[5] = 131;
sin_rom[6] = 157;
sin_rom[7] = 184;
sin_rom[8] = 210;
sin_rom[9] = 236;
sin_rom[10] = 263;
sin_rom[11] = 289;
sin_rom[12] = 315;
sin_rom[13] = 342;
sin_rom[14] = 368;
sin_rom[15] = 394;
sin_rom[16] = 421;
sin_rom[17] = 447;
sin_rom[18] = 473;
sin_rom[19] = 499;
sin_rom[20] = 526;
sin_rom[21] = 552;
sin_rom[22] = 578;
sin_rom[23] = 605;
sin_rom[24] = 631;
sin_rom[25] = 657;
sin_rom[26] = 683;
sin_rom[27] = 709;
sin_rom[28] = 736;
sin_rom[29] = 762;
sin_rom[30] = 788;
sin_rom[31] = 814;
sin_rom[32] = 841;
sin_rom[33] = 867;
sin_rom[34] = 893;
sin_rom[35] = 919;
sin_rom[36] = 945;
sin_rom[37] = 971;
sin_rom[38] = 997;
sin_rom[39] = 1024;
sin_rom[40] = 1050;
sin_rom[41] = 1076;
sin_rom[42] = 1102;
sin_rom[43] = 1128;
sin_rom[44] = 1154;
sin_rom[45] = 1180;
sin_rom[46] = 1206;
sin_rom[47] = 1232;
sin_rom[48] = 1258;
sin_rom[49] = 1284;
sin_rom[50] = 1310;
sin_rom[51] = 1336;
sin_rom[52] = 1362;
sin_rom[53] = 1388;
sin_rom[54] = 1414;
sin_rom[55] = 1440;
sin_rom[56] = 1466;
sin_rom[57] = 1492;
sin_rom[58] = 1518;
sin_rom[59] = 1544;
sin_rom[60] = 1569;
sin_rom[61] = 1595;
sin_rom[62] = 1621;
sin_rom[63] = 1647;
sin_rom[64] = 1673;
sin_rom[65] = 1698;
sin_rom[66] = 1724;
sin_rom[67] = 1750;
sin_rom[68] = 1776;
sin_rom[69] = 1801;
sin_rom[70] = 1827;
sin_rom[71] = 1853;
sin_rom[72] = 1878;
sin_rom[73] = 1904;
sin_rom[74] = 1929;
sin_rom[75] = 1955;
sin_rom[76] = 1981;
sin_rom[77] = 2006;
sin_rom[78] = 2032;
sin_rom[79] = 2057;
sin_rom[80] = 2083;
sin_rom[81] = 2108;
sin_rom[82] = 2134;
sin_rom[83] = 2159;
sin_rom[84] = 2184;
sin_rom[85] = 2210;
sin_rom[86] = 2235;
sin_rom[87] = 2260;
sin_rom[88] = 2286;
sin_rom[89] = 2311;
sin_rom[90] = 2336;
sin_rom[91] = 2361;
sin_rom[92] = 2387;
sin_rom[93] = 2412;
sin_rom[94] = 2437;
sin_rom[95] = 2462;
sin_rom[96] = 2487;
sin_rom[97] = 2512;
sin_rom[98] = 2537;
sin_rom[99] = 2562;
sin_rom[100] = 2587;
sin_rom[101] = 2612;
sin_rom[102] = 2637;
sin_rom[103] = 2662;
sin_rom[104] = 2687;
sin_rom[105] = 2712;
sin_rom[106] = 2737;
sin_rom[107] = 2761;
sin_rom[108] = 2786;
sin_rom[109] = 2811;
sin_rom[110] = 2836;
sin_rom[111] = 2860;
sin_rom[112] = 2885;
sin_rom[113] = 2910;
sin_rom[114] = 2934;
sin_rom[115] = 2959;
sin_rom[116] = 2983;
sin_rom[117] = 3008;
sin_rom[118] = 3032;
sin_rom[119] = 3057;
sin_rom[120] = 3081;
sin_rom[121] = 3106;
sin_rom[122] = 3130;
sin_rom[123] = 3154;
sin_rom[124] = 3178;
sin_rom[125] = 3203;
sin_rom[126] = 3227;
sin_rom[127] = 3251;
sin_rom[128] = 3275;
sin_rom[129] = 3299;
sin_rom[130] = 3323;
sin_rom[131] = 3348;
sin_rom[132] = 3372;
sin_rom[133] = 3396;
sin_rom[134] = 3419;
sin_rom[135] = 3443;
sin_rom[136] = 3467;
sin_rom[137] = 3491;
sin_rom[138] = 3515;
sin_rom[139] = 3539;
sin_rom[140] = 3562;
sin_rom[141] = 3586;
sin_rom[142] = 3610;
sin_rom[143] = 3633;
sin_rom[144] = 3657;
sin_rom[145] = 3680;
sin_rom[146] = 3704;
sin_rom[147] = 3727;
sin_rom[148] = 3751;
sin_rom[149] = 3774;
sin_rom[150] = 3798;
sin_rom[151] = 3821;
sin_rom[152] = 3844;
sin_rom[153] = 3867;
sin_rom[154] = 3891;
sin_rom[155] = 3914;
sin_rom[156] = 3937;
sin_rom[157] = 3960;
sin_rom[158] = 3983;
sin_rom[159] = 4006;
sin_rom[160] = 4029;
sin_rom[161] = 4052;
sin_rom[162] = 4075;
sin_rom[163] = 4097;
sin_rom[164] = 4120;
sin_rom[165] = 4143;
sin_rom[166] = 4166;
sin_rom[167] = 4188;
sin_rom[168] = 4211;
sin_rom[169] = 4233;
sin_rom[170] = 4256;
sin_rom[171] = 4278;
sin_rom[172] = 4301;
sin_rom[173] = 4323;
sin_rom[174] = 4346;
sin_rom[175] = 4368;
sin_rom[176] = 4390;
sin_rom[177] = 4412;
sin_rom[178] = 4434;
sin_rom[179] = 4457;
sin_rom[180] = 4479;
sin_rom[181] = 4501;
sin_rom[182] = 4523;
sin_rom[183] = 4545;
sin_rom[184] = 4566;
sin_rom[185] = 4588;
sin_rom[186] = 4610;
sin_rom[187] = 4632;
sin_rom[188] = 4654;
sin_rom[189] = 4675;
sin_rom[190] = 4697;
sin_rom[191] = 4718;
sin_rom[192] = 4740;
sin_rom[193] = 4761;
sin_rom[194] = 4783;
sin_rom[195] = 4804;
sin_rom[196] = 4825;
sin_rom[197] = 4847;
sin_rom[198] = 4868;
sin_rom[199] = 4889;
sin_rom[200] = 4910;
sin_rom[201] = 4931;
sin_rom[202] = 4952;
sin_rom[203] = 4973;
sin_rom[204] = 4994;
sin_rom[205] = 5015;
sin_rom[206] = 5036;
sin_rom[207] = 5056;
sin_rom[208] = 5077;
sin_rom[209] = 5098;
sin_rom[210] = 5118;
sin_rom[211] = 5139;
sin_rom[212] = 5159;
sin_rom[213] = 5180;
sin_rom[214] = 5200;
sin_rom[215] = 5220;
sin_rom[216] = 5241;
sin_rom[217] = 5261;
sin_rom[218] = 5281;
sin_rom[219] = 5301;
sin_rom[220] = 5321;
sin_rom[221] = 5341;
sin_rom[222] = 5361;
sin_rom[223] = 5381;
sin_rom[224] = 5401;
sin_rom[225] = 5420;
sin_rom[226] = 5440;
sin_rom[227] = 5460;
sin_rom[228] = 5479;
sin_rom[229] = 5499;
sin_rom[230] = 5518;
sin_rom[231] = 5538;
sin_rom[232] = 5557;
sin_rom[233] = 5577;
sin_rom[234] = 5596;
sin_rom[235] = 5615;
sin_rom[236] = 5634;
sin_rom[237] = 5653;
sin_rom[238] = 5672;
sin_rom[239] = 5691;
sin_rom[240] = 5710;
sin_rom[241] = 5729;
sin_rom[242] = 5748;
sin_rom[243] = 5766;
sin_rom[244] = 5785;
sin_rom[245] = 5804;
sin_rom[246] = 5822;
sin_rom[247] = 5841;
sin_rom[248] = 5859;
sin_rom[249] = 5878;
sin_rom[250] = 5896;
sin_rom[251] = 5914;
sin_rom[252] = 5932;
sin_rom[253] = 5950;
sin_rom[254] = 5969;
sin_rom[255] = 5987;
sin_rom[256] = 6004;
sin_rom[257] = 6022;
sin_rom[258] = 6040;
sin_rom[259] = 6058;
sin_rom[260] = 6076;
sin_rom[261] = 6093;
sin_rom[262] = 6111;
sin_rom[263] = 6128;
sin_rom[264] = 6146;
sin_rom[265] = 6163;
sin_rom[266] = 6180;
sin_rom[267] = 6198;
sin_rom[268] = 6215;
sin_rom[269] = 6232;
sin_rom[270] = 6249;
sin_rom[271] = 6266;
sin_rom[272] = 6283;
sin_rom[273] = 6300;
sin_rom[274] = 6317;
sin_rom[275] = 6333;
sin_rom[276] = 6350;
sin_rom[277] = 6367;
sin_rom[278] = 6383;
sin_rom[279] = 6400;
sin_rom[280] = 6416;
sin_rom[281] = 6432;
sin_rom[282] = 6449;
sin_rom[283] = 6465;
sin_rom[284] = 6481;
sin_rom[285] = 6497;
sin_rom[286] = 6513;
sin_rom[287] = 6529;
sin_rom[288] = 6545;
sin_rom[289] = 6561;
sin_rom[290] = 6576;
sin_rom[291] = 6592;
sin_rom[292] = 6608;
sin_rom[293] = 6623;
sin_rom[294] = 6639;
sin_rom[295] = 6654;
sin_rom[296] = 6669;
sin_rom[297] = 6685;
sin_rom[298] = 6700;
sin_rom[299] = 6715;
sin_rom[300] = 6730;
sin_rom[301] = 6745;
sin_rom[302] = 6760;
sin_rom[303] = 6775;
sin_rom[304] = 6789;
sin_rom[305] = 6804;
sin_rom[306] = 6819;
sin_rom[307] = 6833;
sin_rom[308] = 6848;
sin_rom[309] = 6862;
sin_rom[310] = 6876;
sin_rom[311] = 6891;
sin_rom[312] = 6905;
sin_rom[313] = 6919;
sin_rom[314] = 6933;
sin_rom[315] = 6947;
sin_rom[316] = 6961;
sin_rom[317] = 6975;
sin_rom[318] = 6989;
sin_rom[319] = 7002;
sin_rom[320] = 7016;
sin_rom[321] = 7030;
sin_rom[322] = 7043;
sin_rom[323] = 7056;
sin_rom[324] = 7070;
sin_rom[325] = 7083;
sin_rom[326] = 7096;
sin_rom[327] = 7109;
sin_rom[328] = 7122;
sin_rom[329] = 7135;
sin_rom[330] = 7148;
sin_rom[331] = 7161;
sin_rom[332] = 7174;
sin_rom[333] = 7186;
sin_rom[334] = 7199;
sin_rom[335] = 7212;
sin_rom[336] = 7224;
sin_rom[337] = 7236;
sin_rom[338] = 7249;
sin_rom[339] = 7261;
sin_rom[340] = 7273;
sin_rom[341] = 7285;
sin_rom[342] = 7297;
sin_rom[343] = 7309;
sin_rom[344] = 7321;
sin_rom[345] = 7333;
sin_rom[346] = 7344;
sin_rom[347] = 7356;
sin_rom[348] = 7368;
sin_rom[349] = 7379;
sin_rom[350] = 7390;
sin_rom[351] = 7402;
sin_rom[352] = 7413;
sin_rom[353] = 7424;
sin_rom[354] = 7435;
sin_rom[355] = 7446;
sin_rom[356] = 7457;
sin_rom[357] = 7468;
sin_rom[358] = 7479;
sin_rom[359] = 7490;
sin_rom[360] = 7500;
sin_rom[361] = 7511;
sin_rom[362] = 7521;
sin_rom[363] = 7532;
sin_rom[364] = 7542;
sin_rom[365] = 7552;
sin_rom[366] = 7562;
sin_rom[367] = 7572;
sin_rom[368] = 7582;
sin_rom[369] = 7592;
sin_rom[370] = 7602;
sin_rom[371] = 7612;
sin_rom[372] = 7622;
sin_rom[373] = 7631;
sin_rom[374] = 7641;
sin_rom[375] = 7650;
sin_rom[376] = 7660;
sin_rom[377] = 7669;
sin_rom[378] = 7678;
sin_rom[379] = 7687;
sin_rom[380] = 7696;
sin_rom[381] = 7705;
sin_rom[382] = 7714;
sin_rom[383] = 7723;
sin_rom[384] = 7732;
sin_rom[385] = 7740;
sin_rom[386] = 7749;
sin_rom[387] = 7757;
sin_rom[388] = 7766;
sin_rom[389] = 7774;
sin_rom[390] = 7782;
sin_rom[391] = 7791;
sin_rom[392] = 7799;
sin_rom[393] = 7807;
sin_rom[394] = 7815;
sin_rom[395] = 7822;
sin_rom[396] = 7830;
sin_rom[397] = 7838;
sin_rom[398] = 7846;
sin_rom[399] = 7853;
sin_rom[400] = 7861;
sin_rom[401] = 7868;
sin_rom[402] = 7875;
sin_rom[403] = 7882;
sin_rom[404] = 7890;
sin_rom[405] = 7897;
sin_rom[406] = 7904;
sin_rom[407] = 7910;
sin_rom[408] = 7917;
sin_rom[409] = 7924;
sin_rom[410] = 7931;
sin_rom[411] = 7937;
sin_rom[412] = 7944;
sin_rom[413] = 7950;
sin_rom[414] = 7956;
sin_rom[415] = 7962;
sin_rom[416] = 7969;
sin_rom[417] = 7975;
sin_rom[418] = 7981;
sin_rom[419] = 7987;
sin_rom[420] = 7992;
sin_rom[421] = 7998;
sin_rom[422] = 8004;
sin_rom[423] = 8009;
sin_rom[424] = 8015;
sin_rom[425] = 8020;
sin_rom[426] = 8025;
sin_rom[427] = 8031;
sin_rom[428] = 8036;
sin_rom[429] = 8041;
sin_rom[430] = 8046;
sin_rom[431] = 8051;
sin_rom[432] = 8056;
sin_rom[433] = 8060;
sin_rom[434] = 8065;
sin_rom[435] = 8070;
sin_rom[436] = 8074;
sin_rom[437] = 8078;
sin_rom[438] = 8083;
sin_rom[439] = 8087;
sin_rom[440] = 8091;
sin_rom[441] = 8095;
sin_rom[442] = 8099;
sin_rom[443] = 8103;
sin_rom[444] = 8107;
sin_rom[445] = 8111;
sin_rom[446] = 8114;
sin_rom[447] = 8118;
sin_rom[448] = 8121;
sin_rom[449] = 8125;
sin_rom[450] = 8128;
sin_rom[451] = 8131;
sin_rom[452] = 8134;
sin_rom[453] = 8137;
sin_rom[454] = 8140;
sin_rom[455] = 8143;
sin_rom[456] = 8146;
sin_rom[457] = 8149;
sin_rom[458] = 8152;
sin_rom[459] = 8154;
sin_rom[460] = 8157;
sin_rom[461] = 8159;
sin_rom[462] = 8161;
sin_rom[463] = 8163;
sin_rom[464] = 8166;
sin_rom[465] = 8168;
sin_rom[466] = 8170;
sin_rom[467] = 8171;
sin_rom[468] = 8173;
sin_rom[469] = 8175;
sin_rom[470] = 8177;
sin_rom[471] = 8178;
sin_rom[472] = 8180;
sin_rom[473] = 8181;
sin_rom[474] = 8182;
sin_rom[475] = 8184;
sin_rom[476] = 8185;
sin_rom[477] = 8186;
sin_rom[478] = 8187;
sin_rom[479] = 8187;
sin_rom[480] = 8188;
sin_rom[481] = 8189;
sin_rom[482] = 8190;
sin_rom[483] = 8190;
sin_rom[484] = 8191;
sin_rom[485] = 8191;
sin_rom[486] = 8191;
sin_rom[487] = 8191;
sin_rom[488] = 8191;
sin_rom[489] = 8191;
sin_rom[490] = 8191;
sin_rom[491] = 8191;
sin_rom[492] = 8191;
sin_rom[493] = 8191;
sin_rom[494] = 8190;
sin_rom[495] = 8190;
sin_rom[496] = 8189;
sin_rom[497] = 8189;
sin_rom[498] = 8188;
sin_rom[499] = 8187;
sin_rom[500] = 8186;
sin_rom[501] = 8185;
sin_rom[502] = 8184;
sin_rom[503] = 8183;
sin_rom[504] = 8182;
sin_rom[505] = 8180;
sin_rom[506] = 8179;
sin_rom[507] = 8177;
sin_rom[508] = 8176;
sin_rom[509] = 8174;
sin_rom[510] = 8172;
sin_rom[511] = 8171;
sin_rom[512] = 8169;
sin_rom[513] = 8167;
sin_rom[514] = 8165;
sin_rom[515] = 8162;
sin_rom[516] = 8160;
sin_rom[517] = 8158;
sin_rom[518] = 8155;
sin_rom[519] = 8153;
sin_rom[520] = 8150;
sin_rom[521] = 8148;
sin_rom[522] = 8145;
sin_rom[523] = 8142;
sin_rom[524] = 8139;
sin_rom[525] = 8136;
sin_rom[526] = 8133;
sin_rom[527] = 8130;
sin_rom[528] = 8126;
sin_rom[529] = 8123;
sin_rom[530] = 8120;
sin_rom[531] = 8116;
sin_rom[532] = 8112;
sin_rom[533] = 8109;
sin_rom[534] = 8105;
sin_rom[535] = 8101;
sin_rom[536] = 8097;
sin_rom[537] = 8093;
sin_rom[538] = 8089;
sin_rom[539] = 8085;
sin_rom[540] = 8081;
sin_rom[541] = 8076;
sin_rom[542] = 8072;
sin_rom[543] = 8067;
sin_rom[544] = 8063;
sin_rom[545] = 8058;
sin_rom[546] = 8053;
sin_rom[547] = 8048;
sin_rom[548] = 8043;
sin_rom[549] = 8038;
sin_rom[550] = 8033;
sin_rom[551] = 8028;
sin_rom[552] = 8023;
sin_rom[553] = 8017;
sin_rom[554] = 8012;
sin_rom[555] = 8006;
sin_rom[556] = 8001;
sin_rom[557] = 7995;
sin_rom[558] = 7989;
sin_rom[559] = 7984;
sin_rom[560] = 7978;
sin_rom[561] = 7972;
sin_rom[562] = 7966;
sin_rom[563] = 7959;
sin_rom[564] = 7953;
sin_rom[565] = 7947;
sin_rom[566] = 7940;
sin_rom[567] = 7934;
sin_rom[568] = 7927;
sin_rom[569] = 7921;
sin_rom[570] = 7914;
sin_rom[571] = 7907;
sin_rom[572] = 7900;
sin_rom[573] = 7893;
sin_rom[574] = 7886;
sin_rom[575] = 7879;
sin_rom[576] = 7872;
sin_rom[577] = 7864;
sin_rom[578] = 7857;
sin_rom[579] = 7849;
sin_rom[580] = 7842;
sin_rom[581] = 7834;
sin_rom[582] = 7826;
sin_rom[583] = 7819;
sin_rom[584] = 7811;
sin_rom[585] = 7803;
sin_rom[586] = 7795;
sin_rom[587] = 7786;
sin_rom[588] = 7778;
sin_rom[589] = 7770;
sin_rom[590] = 7762;
sin_rom[591] = 7753;
sin_rom[592] = 7745;
sin_rom[593] = 7736;
sin_rom[594] = 7727;
sin_rom[595] = 7718;
sin_rom[596] = 7710;
sin_rom[597] = 7701;
sin_rom[598] = 7692;
sin_rom[599] = 7683;
sin_rom[600] = 7673;
sin_rom[601] = 7664;
sin_rom[602] = 7655;
sin_rom[603] = 7645;
sin_rom[604] = 7636;
sin_rom[605] = 7626;
sin_rom[606] = 7617;
sin_rom[607] = 7607;
sin_rom[608] = 7597;
sin_rom[609] = 7587;
sin_rom[610] = 7577;
sin_rom[611] = 7567;
sin_rom[612] = 7557;
sin_rom[613] = 7547;
sin_rom[614] = 7537;
sin_rom[615] = 7526;
sin_rom[616] = 7516;
sin_rom[617] = 7505;
sin_rom[618] = 7495;
sin_rom[619] = 7484;
sin_rom[620] = 7473;
sin_rom[621] = 7463;
sin_rom[622] = 7452;
sin_rom[623] = 7441;
sin_rom[624] = 7430;
sin_rom[625] = 7419;
sin_rom[626] = 7407;
sin_rom[627] = 7396;
sin_rom[628] = 7385;
sin_rom[629] = 7373;
sin_rom[630] = 7362;
sin_rom[631] = 7350;
sin_rom[632] = 7339;
sin_rom[633] = 7327;
sin_rom[634] = 7315;
sin_rom[635] = 7303;
sin_rom[636] = 7291;
sin_rom[637] = 7279;
sin_rom[638] = 7267;
sin_rom[639] = 7255;
sin_rom[640] = 7243;
sin_rom[641] = 7230;
sin_rom[642] = 7218;
sin_rom[643] = 7205;
sin_rom[644] = 7193;
sin_rom[645] = 7180;
sin_rom[646] = 7167;
sin_rom[647] = 7155;
sin_rom[648] = 7142;
sin_rom[649] = 7129;
sin_rom[650] = 7116;
sin_rom[651] = 7103;
sin_rom[652] = 7090;
sin_rom[653] = 7076;
sin_rom[654] = 7063;
sin_rom[655] = 7050;
sin_rom[656] = 7036;
sin_rom[657] = 7023;
sin_rom[658] = 7009;
sin_rom[659] = 6995;
sin_rom[660] = 6982;
sin_rom[661] = 6968;
sin_rom[662] = 6954;
sin_rom[663] = 6940;
sin_rom[664] = 6926;
sin_rom[665] = 6912;
sin_rom[666] = 6898;
sin_rom[667] = 6884;
sin_rom[668] = 6869;
sin_rom[669] = 6855;
sin_rom[670] = 6840;
sin_rom[671] = 6826;
sin_rom[672] = 6811;
sin_rom[673] = 6797;
sin_rom[674] = 6782;
sin_rom[675] = 6767;
sin_rom[676] = 6752;
sin_rom[677] = 6737;
sin_rom[678] = 6722;
sin_rom[679] = 6707;
sin_rom[680] = 6692;
sin_rom[681] = 6677;
sin_rom[682] = 6662;
sin_rom[683] = 6646;
sin_rom[684] = 6631;
sin_rom[685] = 6615;
sin_rom[686] = 6600;
sin_rom[687] = 6584;
sin_rom[688] = 6568;
sin_rom[689] = 6553;
sin_rom[690] = 6537;
sin_rom[691] = 6521;
sin_rom[692] = 6505;
sin_rom[693] = 6489;
sin_rom[694] = 6473;
sin_rom[695] = 6457;
sin_rom[696] = 6440;
sin_rom[697] = 6424;
sin_rom[698] = 6408;
sin_rom[699] = 6391;
sin_rom[700] = 6375;
sin_rom[701] = 6358;
sin_rom[702] = 6342;
sin_rom[703] = 6325;
sin_rom[704] = 6308;
sin_rom[705] = 6291;
sin_rom[706] = 6274;
sin_rom[707] = 6257;
sin_rom[708] = 6240;
sin_rom[709] = 6223;
sin_rom[710] = 6206;
sin_rom[711] = 6189;
sin_rom[712] = 6172;
sin_rom[713] = 6154;
sin_rom[714] = 6137;
sin_rom[715] = 6119;
sin_rom[716] = 6102;
sin_rom[717] = 6084;
sin_rom[718] = 6067;
sin_rom[719] = 6049;
sin_rom[720] = 6031;
sin_rom[721] = 6013;
sin_rom[722] = 5995;
sin_rom[723] = 5977;
sin_rom[724] = 5959;
sin_rom[725] = 5941;
sin_rom[726] = 5923;
sin_rom[727] = 5905;
sin_rom[728] = 5887;
sin_rom[729] = 5868;
sin_rom[730] = 5850;
sin_rom[731] = 5831;
sin_rom[732] = 5813;
sin_rom[733] = 5794;
sin_rom[734] = 5776;
sin_rom[735] = 5757;
sin_rom[736] = 5738;
sin_rom[737] = 5719;
sin_rom[738] = 5701;
sin_rom[739] = 5682;
sin_rom[740] = 5663;
sin_rom[741] = 5644;
sin_rom[742] = 5624;
sin_rom[743] = 5605;
sin_rom[744] = 5586;
sin_rom[745] = 5567;
sin_rom[746] = 5547;
sin_rom[747] = 5528;
sin_rom[748] = 5509;
sin_rom[749] = 5489;
sin_rom[750] = 5470;
sin_rom[751] = 5450;
sin_rom[752] = 5430;
sin_rom[753] = 5410;
sin_rom[754] = 5391;
sin_rom[755] = 5371;
sin_rom[756] = 5351;
sin_rom[757] = 5331;
sin_rom[758] = 5311;
sin_rom[759] = 5291;
sin_rom[760] = 5271;
sin_rom[761] = 5251;
sin_rom[762] = 5230;
sin_rom[763] = 5210;
sin_rom[764] = 5190;
sin_rom[765] = 5169;
sin_rom[766] = 5149;
sin_rom[767] = 5128;
sin_rom[768] = 5108;
sin_rom[769] = 5087;
sin_rom[770] = 5067;
sin_rom[771] = 5046;
sin_rom[772] = 5025;
sin_rom[773] = 5004;
sin_rom[774] = 4983;
sin_rom[775] = 4962;
sin_rom[776] = 4941;
sin_rom[777] = 4920;
sin_rom[778] = 4899;
sin_rom[779] = 4878;
sin_rom[780] = 4857;
sin_rom[781] = 4836;
sin_rom[782] = 4815;
sin_rom[783] = 4793;
sin_rom[784] = 4772;
sin_rom[785] = 4750;
sin_rom[786] = 4729;
sin_rom[787] = 4707;
sin_rom[788] = 4686;
sin_rom[789] = 4664;
sin_rom[790] = 4643;
sin_rom[791] = 4621;
sin_rom[792] = 4599;
sin_rom[793] = 4577;
sin_rom[794] = 4555;
sin_rom[795] = 4534;
sin_rom[796] = 4512;
sin_rom[797] = 4490;
sin_rom[798] = 4468;
sin_rom[799] = 4445;
sin_rom[800] = 4423;
sin_rom[801] = 4401;
sin_rom[802] = 4379;
sin_rom[803] = 4357;
sin_rom[804] = 4334;
sin_rom[805] = 4312;
sin_rom[806] = 4290;
sin_rom[807] = 4267;
sin_rom[808] = 4245;
sin_rom[809] = 4222;
sin_rom[810] = 4199;
sin_rom[811] = 4177;
sin_rom[812] = 4154;
sin_rom[813] = 4131;
sin_rom[814] = 4109;
sin_rom[815] = 4086;
sin_rom[816] = 4063;
sin_rom[817] = 4040;
sin_rom[818] = 4017;
sin_rom[819] = 3994;
sin_rom[820] = 3971;
sin_rom[821] = 3948;
sin_rom[822] = 3925;
sin_rom[823] = 3902;
sin_rom[824] = 3879;
sin_rom[825] = 3856;
sin_rom[826] = 3832;
sin_rom[827] = 3809;
sin_rom[828] = 3786;
sin_rom[829] = 3762;
sin_rom[830] = 3739;
sin_rom[831] = 3716;
sin_rom[832] = 3692;
sin_rom[833] = 3669;
sin_rom[834] = 3645;
sin_rom[835] = 3621;
sin_rom[836] = 3598;
sin_rom[837] = 3574;
sin_rom[838] = 3550;
sin_rom[839] = 3527;
sin_rom[840] = 3503;
sin_rom[841] = 3479;
sin_rom[842] = 3455;
sin_rom[843] = 3431;
sin_rom[844] = 3407;
sin_rom[845] = 3383;
sin_rom[846] = 3359;
sin_rom[847] = 3335;
sin_rom[848] = 3311;
sin_rom[849] = 3287;
sin_rom[850] = 3263;
sin_rom[851] = 3239;
sin_rom[852] = 3215;
sin_rom[853] = 3191;
sin_rom[854] = 3166;
sin_rom[855] = 3142;
sin_rom[856] = 3118;
sin_rom[857] = 3093;
sin_rom[858] = 3069;
sin_rom[859] = 3044;
sin_rom[860] = 3020;
sin_rom[861] = 2995;
sin_rom[862] = 2971;
sin_rom[863] = 2946;
sin_rom[864] = 2922;
sin_rom[865] = 2897;
sin_rom[866] = 2873;
sin_rom[867] = 2848;
sin_rom[868] = 2823;
sin_rom[869] = 2798;
sin_rom[870] = 2774;
sin_rom[871] = 2749;
sin_rom[872] = 2724;
sin_rom[873] = 2699;
sin_rom[874] = 2674;
sin_rom[875] = 2650;
sin_rom[876] = 2625;
sin_rom[877] = 2600;
sin_rom[878] = 2575;
sin_rom[879] = 2550;
sin_rom[880] = 2525;
sin_rom[881] = 2500;
sin_rom[882] = 2474;
sin_rom[883] = 2449;
sin_rom[884] = 2424;
sin_rom[885] = 2399;
sin_rom[886] = 2374;
sin_rom[887] = 2349;
sin_rom[888] = 2323;
sin_rom[889] = 2298;
sin_rom[890] = 2273;
sin_rom[891] = 2248;
sin_rom[892] = 2222;
sin_rom[893] = 2197;
sin_rom[894] = 2172;
sin_rom[895] = 2146;
sin_rom[896] = 2121;
sin_rom[897] = 2095;
sin_rom[898] = 2070;
sin_rom[899] = 2044;
sin_rom[900] = 2019;
sin_rom[901] = 1993;
sin_rom[902] = 1968;
sin_rom[903] = 1942;
sin_rom[904] = 1917;
sin_rom[905] = 1891;
sin_rom[906] = 1865;
sin_rom[907] = 1840;
sin_rom[908] = 1814;
sin_rom[909] = 1788;
sin_rom[910] = 1763;
sin_rom[911] = 1737;
sin_rom[912] = 1711;
sin_rom[913] = 1685;
sin_rom[914] = 1660;
sin_rom[915] = 1634;
sin_rom[916] = 1608;
sin_rom[917] = 1582;
sin_rom[918] = 1556;
sin_rom[919] = 1531;
sin_rom[920] = 1505;
sin_rom[921] = 1479;
sin_rom[922] = 1453;
sin_rom[923] = 1427;
sin_rom[924] = 1401;
sin_rom[925] = 1375;
sin_rom[926] = 1349;
sin_rom[927] = 1323;
sin_rom[928] = 1297;
sin_rom[929] = 1271;
sin_rom[930] = 1245;
sin_rom[931] = 1219;
sin_rom[932] = 1193;
sin_rom[933] = 1167;
sin_rom[934] = 1141;
sin_rom[935] = 1115;
sin_rom[936] = 1089;
sin_rom[937] = 1063;
sin_rom[938] = 1037;
sin_rom[939] = 1010;
sin_rom[940] = 984;
sin_rom[941] = 958;
sin_rom[942] = 932;
sin_rom[943] = 906;
sin_rom[944] = 880;
sin_rom[945] = 854;
sin_rom[946] = 827;
sin_rom[947] = 801;
sin_rom[948] = 775;
sin_rom[949] = 749;
sin_rom[950] = 722;
sin_rom[951] = 696;
sin_rom[952] = 670;
sin_rom[953] = 644;
sin_rom[954] = 618;
sin_rom[955] = 591;
sin_rom[956] = 565;
sin_rom[957] = 539;
sin_rom[958] = 512;
sin_rom[959] = 486;
sin_rom[960] = 460;
sin_rom[961] = 434;
sin_rom[962] = 407;
sin_rom[963] = 381;
sin_rom[964] = 355;
sin_rom[965] = 328;
sin_rom[966] = 302;
sin_rom[967] = 276;
sin_rom[968] = 249;
sin_rom[969] = 223;
sin_rom[970] = 197;
sin_rom[971] = 171;
sin_rom[972] = 144;
sin_rom[973] = 118;
sin_rom[974] = 92;
sin_rom[975] = 65;
sin_rom[976] = 39;
sin_rom[977] = 13;
sin_rom[978] = -13;
sin_rom[979] = -39;
sin_rom[980] = -65;
sin_rom[981] = -92;
sin_rom[982] = -118;
sin_rom[983] = -144;
sin_rom[984] = -171;
sin_rom[985] = -197;
sin_rom[986] = -223;
sin_rom[987] = -250;
sin_rom[988] = -276;
sin_rom[989] = -302;
sin_rom[990] = -329;
sin_rom[991] = -355;
sin_rom[992] = -381;
sin_rom[993] = -408;
sin_rom[994] = -434;
sin_rom[995] = -460;
sin_rom[996] = -486;
sin_rom[997] = -513;
sin_rom[998] = -539;
sin_rom[999] = -565;
sin_rom[1000] = -591;
sin_rom[1001] = -618;
sin_rom[1002] = -644;
sin_rom[1003] = -670;
sin_rom[1004] = -696;
sin_rom[1005] = -723;
sin_rom[1006] = -749;
sin_rom[1007] = -775;
sin_rom[1008] = -801;
sin_rom[1009] = -828;
sin_rom[1010] = -854;
sin_rom[1011] = -880;
sin_rom[1012] = -906;
sin_rom[1013] = -932;
sin_rom[1014] = -958;
sin_rom[1015] = -985;
sin_rom[1016] = -1011;
sin_rom[1017] = -1037;
sin_rom[1018] = -1063;
sin_rom[1019] = -1089;
sin_rom[1020] = -1115;
sin_rom[1021] = -1141;
sin_rom[1022] = -1167;
sin_rom[1023] = -1193;
sin_rom[1024] = -1219;
sin_rom[1025] = -1245;
sin_rom[1026] = -1271;
sin_rom[1027] = -1297;
sin_rom[1028] = -1323;
sin_rom[1029] = -1349;
sin_rom[1030] = -1375;
sin_rom[1031] = -1401;
sin_rom[1032] = -1427;
sin_rom[1033] = -1453;
sin_rom[1034] = -1479;
sin_rom[1035] = -1505;
sin_rom[1036] = -1531;
sin_rom[1037] = -1557;
sin_rom[1038] = -1582;
sin_rom[1039] = -1608;
sin_rom[1040] = -1634;
sin_rom[1041] = -1660;
sin_rom[1042] = -1686;
sin_rom[1043] = -1711;
sin_rom[1044] = -1737;
sin_rom[1045] = -1763;
sin_rom[1046] = -1789;
sin_rom[1047] = -1814;
sin_rom[1048] = -1840;
sin_rom[1049] = -1866;
sin_rom[1050] = -1891;
sin_rom[1051] = -1917;
sin_rom[1052] = -1942;
sin_rom[1053] = -1968;
sin_rom[1054] = -1994;
sin_rom[1055] = -2019;
sin_rom[1056] = -2045;
sin_rom[1057] = -2070;
sin_rom[1058] = -2095;
sin_rom[1059] = -2121;
sin_rom[1060] = -2146;
sin_rom[1061] = -2172;
sin_rom[1062] = -2197;
sin_rom[1063] = -2222;
sin_rom[1064] = -2248;
sin_rom[1065] = -2273;
sin_rom[1066] = -2298;
sin_rom[1067] = -2324;
sin_rom[1068] = -2349;
sin_rom[1069] = -2374;
sin_rom[1070] = -2399;
sin_rom[1071] = -2424;
sin_rom[1072] = -2450;
sin_rom[1073] = -2475;
sin_rom[1074] = -2500;
sin_rom[1075] = -2525;
sin_rom[1076] = -2550;
sin_rom[1077] = -2575;
sin_rom[1078] = -2600;
sin_rom[1079] = -2625;
sin_rom[1080] = -2650;
sin_rom[1081] = -2675;
sin_rom[1082] = -2699;
sin_rom[1083] = -2724;
sin_rom[1084] = -2749;
sin_rom[1085] = -2774;
sin_rom[1086] = -2799;
sin_rom[1087] = -2823;
sin_rom[1088] = -2848;
sin_rom[1089] = -2873;
sin_rom[1090] = -2897;
sin_rom[1091] = -2922;
sin_rom[1092] = -2947;
sin_rom[1093] = -2971;
sin_rom[1094] = -2996;
sin_rom[1095] = -3020;
sin_rom[1096] = -3045;
sin_rom[1097] = -3069;
sin_rom[1098] = -3093;
sin_rom[1099] = -3118;
sin_rom[1100] = -3142;
sin_rom[1101] = -3166;
sin_rom[1102] = -3191;
sin_rom[1103] = -3215;
sin_rom[1104] = -3239;
sin_rom[1105] = -3263;
sin_rom[1106] = -3287;
sin_rom[1107] = -3312;
sin_rom[1108] = -3336;
sin_rom[1109] = -3360;
sin_rom[1110] = -3384;
sin_rom[1111] = -3408;
sin_rom[1112] = -3432;
sin_rom[1113] = -3455;
sin_rom[1114] = -3479;
sin_rom[1115] = -3503;
sin_rom[1116] = -3527;
sin_rom[1117] = -3551;
sin_rom[1118] = -3574;
sin_rom[1119] = -3598;
sin_rom[1120] = -3622;
sin_rom[1121] = -3645;
sin_rom[1122] = -3669;
sin_rom[1123] = -3692;
sin_rom[1124] = -3716;
sin_rom[1125] = -3739;
sin_rom[1126] = -3763;
sin_rom[1127] = -3786;
sin_rom[1128] = -3809;
sin_rom[1129] = -3833;
sin_rom[1130] = -3856;
sin_rom[1131] = -3879;
sin_rom[1132] = -3902;
sin_rom[1133] = -3925;
sin_rom[1134] = -3948;
sin_rom[1135] = -3971;
sin_rom[1136] = -3995;
sin_rom[1137] = -4017;
sin_rom[1138] = -4040;
sin_rom[1139] = -4063;
sin_rom[1140] = -4086;
sin_rom[1141] = -4109;
sin_rom[1142] = -4132;
sin_rom[1143] = -4154;
sin_rom[1144] = -4177;
sin_rom[1145] = -4200;
sin_rom[1146] = -4222;
sin_rom[1147] = -4245;
sin_rom[1148] = -4267;
sin_rom[1149] = -4290;
sin_rom[1150] = -4312;
sin_rom[1151] = -4335;
sin_rom[1152] = -4357;
sin_rom[1153] = -4379;
sin_rom[1154] = -4401;
sin_rom[1155] = -4424;
sin_rom[1156] = -4446;
sin_rom[1157] = -4468;
sin_rom[1158] = -4490;
sin_rom[1159] = -4512;
sin_rom[1160] = -4534;
sin_rom[1161] = -4556;
sin_rom[1162] = -4577;
sin_rom[1163] = -4599;
sin_rom[1164] = -4621;
sin_rom[1165] = -4643;
sin_rom[1166] = -4664;
sin_rom[1167] = -4686;
sin_rom[1168] = -4708;
sin_rom[1169] = -4729;
sin_rom[1170] = -4751;
sin_rom[1171] = -4772;
sin_rom[1172] = -4793;
sin_rom[1173] = -4815;
sin_rom[1174] = -4836;
sin_rom[1175] = -4857;
sin_rom[1176] = -4878;
sin_rom[1177] = -4900;
sin_rom[1178] = -4921;
sin_rom[1179] = -4942;
sin_rom[1180] = -4963;
sin_rom[1181] = -4984;
sin_rom[1182] = -5004;
sin_rom[1183] = -5025;
sin_rom[1184] = -5046;
sin_rom[1185] = -5067;
sin_rom[1186] = -5087;
sin_rom[1187] = -5108;
sin_rom[1188] = -5129;
sin_rom[1189] = -5149;
sin_rom[1190] = -5169;
sin_rom[1191] = -5190;
sin_rom[1192] = -5210;
sin_rom[1193] = -5231;
sin_rom[1194] = -5251;
sin_rom[1195] = -5271;
sin_rom[1196] = -5291;
sin_rom[1197] = -5311;
sin_rom[1198] = -5331;
sin_rom[1199] = -5351;
sin_rom[1200] = -5371;
sin_rom[1201] = -5391;
sin_rom[1202] = -5411;
sin_rom[1203] = -5430;
sin_rom[1204] = -5450;
sin_rom[1205] = -5470;
sin_rom[1206] = -5489;
sin_rom[1207] = -5509;
sin_rom[1208] = -5528;
sin_rom[1209] = -5548;
sin_rom[1210] = -5567;
sin_rom[1211] = -5586;
sin_rom[1212] = -5605;
sin_rom[1213] = -5625;
sin_rom[1214] = -5644;
sin_rom[1215] = -5663;
sin_rom[1216] = -5682;
sin_rom[1217] = -5701;
sin_rom[1218] = -5720;
sin_rom[1219] = -5738;
sin_rom[1220] = -5757;
sin_rom[1221] = -5776;
sin_rom[1222] = -5795;
sin_rom[1223] = -5813;
sin_rom[1224] = -5832;
sin_rom[1225] = -5850;
sin_rom[1226] = -5869;
sin_rom[1227] = -5887;
sin_rom[1228] = -5905;
sin_rom[1229] = -5923;
sin_rom[1230] = -5941;
sin_rom[1231] = -5960;
sin_rom[1232] = -5978;
sin_rom[1233] = -5996;
sin_rom[1234] = -6013;
sin_rom[1235] = -6031;
sin_rom[1236] = -6049;
sin_rom[1237] = -6067;
sin_rom[1238] = -6085;
sin_rom[1239] = -6102;
sin_rom[1240] = -6120;
sin_rom[1241] = -6137;
sin_rom[1242] = -6155;
sin_rom[1243] = -6172;
sin_rom[1244] = -6189;
sin_rom[1245] = -6206;
sin_rom[1246] = -6223;
sin_rom[1247] = -6241;
sin_rom[1248] = -6258;
sin_rom[1249] = -6275;
sin_rom[1250] = -6291;
sin_rom[1251] = -6308;
sin_rom[1252] = -6325;
sin_rom[1253] = -6342;
sin_rom[1254] = -6358;
sin_rom[1255] = -6375;
sin_rom[1256] = -6391;
sin_rom[1257] = -6408;
sin_rom[1258] = -6424;
sin_rom[1259] = -6441;
sin_rom[1260] = -6457;
sin_rom[1261] = -6473;
sin_rom[1262] = -6489;
sin_rom[1263] = -6505;
sin_rom[1264] = -6521;
sin_rom[1265] = -6537;
sin_rom[1266] = -6553;
sin_rom[1267] = -6569;
sin_rom[1268] = -6584;
sin_rom[1269] = -6600;
sin_rom[1270] = -6615;
sin_rom[1271] = -6631;
sin_rom[1272] = -6646;
sin_rom[1273] = -6662;
sin_rom[1274] = -6677;
sin_rom[1275] = -6692;
sin_rom[1276] = -6707;
sin_rom[1277] = -6722;
sin_rom[1278] = -6737;
sin_rom[1279] = -6752;
sin_rom[1280] = -6767;
sin_rom[1281] = -6782;
sin_rom[1282] = -6797;
sin_rom[1283] = -6811;
sin_rom[1284] = -6826;
sin_rom[1285] = -6841;
sin_rom[1286] = -6855;
sin_rom[1287] = -6869;
sin_rom[1288] = -6884;
sin_rom[1289] = -6898;
sin_rom[1290] = -6912;
sin_rom[1291] = -6926;
sin_rom[1292] = -6940;
sin_rom[1293] = -6954;
sin_rom[1294] = -6968;
sin_rom[1295] = -6982;
sin_rom[1296] = -6996;
sin_rom[1297] = -7009;
sin_rom[1298] = -7023;
sin_rom[1299] = -7036;
sin_rom[1300] = -7050;
sin_rom[1301] = -7063;
sin_rom[1302] = -7076;
sin_rom[1303] = -7090;
sin_rom[1304] = -7103;
sin_rom[1305] = -7116;
sin_rom[1306] = -7129;
sin_rom[1307] = -7142;
sin_rom[1308] = -7155;
sin_rom[1309] = -7167;
sin_rom[1310] = -7180;
sin_rom[1311] = -7193;
sin_rom[1312] = -7205;
sin_rom[1313] = -7218;
sin_rom[1314] = -7230;
sin_rom[1315] = -7243;
sin_rom[1316] = -7255;
sin_rom[1317] = -7267;
sin_rom[1318] = -7279;
sin_rom[1319] = -7291;
sin_rom[1320] = -7303;
sin_rom[1321] = -7315;
sin_rom[1322] = -7327;
sin_rom[1323] = -7339;
sin_rom[1324] = -7350;
sin_rom[1325] = -7362;
sin_rom[1326] = -7373;
sin_rom[1327] = -7385;
sin_rom[1328] = -7396;
sin_rom[1329] = -7407;
sin_rom[1330] = -7419;
sin_rom[1331] = -7430;
sin_rom[1332] = -7441;
sin_rom[1333] = -7452;
sin_rom[1334] = -7463;
sin_rom[1335] = -7473;
sin_rom[1336] = -7484;
sin_rom[1337] = -7495;
sin_rom[1338] = -7505;
sin_rom[1339] = -7516;
sin_rom[1340] = -7526;
sin_rom[1341] = -7537;
sin_rom[1342] = -7547;
sin_rom[1343] = -7557;
sin_rom[1344] = -7567;
sin_rom[1345] = -7577;
sin_rom[1346] = -7587;
sin_rom[1347] = -7597;
sin_rom[1348] = -7607;
sin_rom[1349] = -7617;
sin_rom[1350] = -7626;
sin_rom[1351] = -7636;
sin_rom[1352] = -7645;
sin_rom[1353] = -7655;
sin_rom[1354] = -7664;
sin_rom[1355] = -7673;
sin_rom[1356] = -7683;
sin_rom[1357] = -7692;
sin_rom[1358] = -7701;
sin_rom[1359] = -7710;
sin_rom[1360] = -7719;
sin_rom[1361] = -7727;
sin_rom[1362] = -7736;
sin_rom[1363] = -7745;
sin_rom[1364] = -7753;
sin_rom[1365] = -7762;
sin_rom[1366] = -7770;
sin_rom[1367] = -7778;
sin_rom[1368] = -7787;
sin_rom[1369] = -7795;
sin_rom[1370] = -7803;
sin_rom[1371] = -7811;
sin_rom[1372] = -7819;
sin_rom[1373] = -7826;
sin_rom[1374] = -7834;
sin_rom[1375] = -7842;
sin_rom[1376] = -7849;
sin_rom[1377] = -7857;
sin_rom[1378] = -7864;
sin_rom[1379] = -7872;
sin_rom[1380] = -7879;
sin_rom[1381] = -7886;
sin_rom[1382] = -7893;
sin_rom[1383] = -7900;
sin_rom[1384] = -7907;
sin_rom[1385] = -7914;
sin_rom[1386] = -7921;
sin_rom[1387] = -7927;
sin_rom[1388] = -7934;
sin_rom[1389] = -7940;
sin_rom[1390] = -7947;
sin_rom[1391] = -7953;
sin_rom[1392] = -7959;
sin_rom[1393] = -7966;
sin_rom[1394] = -7972;
sin_rom[1395] = -7978;
sin_rom[1396] = -7984;
sin_rom[1397] = -7989;
sin_rom[1398] = -7995;
sin_rom[1399] = -8001;
sin_rom[1400] = -8007;
sin_rom[1401] = -8012;
sin_rom[1402] = -8018;
sin_rom[1403] = -8023;
sin_rom[1404] = -8028;
sin_rom[1405] = -8033;
sin_rom[1406] = -8038;
sin_rom[1407] = -8043;
sin_rom[1408] = -8048;
sin_rom[1409] = -8053;
sin_rom[1410] = -8058;
sin_rom[1411] = -8063;
sin_rom[1412] = -8067;
sin_rom[1413] = -8072;
sin_rom[1414] = -8076;
sin_rom[1415] = -8081;
sin_rom[1416] = -8085;
sin_rom[1417] = -8089;
sin_rom[1418] = -8093;
sin_rom[1419] = -8097;
sin_rom[1420] = -8101;
sin_rom[1421] = -8105;
sin_rom[1422] = -8109;
sin_rom[1423] = -8113;
sin_rom[1424] = -8116;
sin_rom[1425] = -8120;
sin_rom[1426] = -8123;
sin_rom[1427] = -8126;
sin_rom[1428] = -8130;
sin_rom[1429] = -8133;
sin_rom[1430] = -8136;
sin_rom[1431] = -8139;
sin_rom[1432] = -8142;
sin_rom[1433] = -8145;
sin_rom[1434] = -8148;
sin_rom[1435] = -8150;
sin_rom[1436] = -8153;
sin_rom[1437] = -8155;
sin_rom[1438] = -8158;
sin_rom[1439] = -8160;
sin_rom[1440] = -8162;
sin_rom[1441] = -8165;
sin_rom[1442] = -8167;
sin_rom[1443] = -8169;
sin_rom[1444] = -8171;
sin_rom[1445] = -8172;
sin_rom[1446] = -8174;
sin_rom[1447] = -8176;
sin_rom[1448] = -8177;
sin_rom[1449] = -8179;
sin_rom[1450] = -8180;
sin_rom[1451] = -8182;
sin_rom[1452] = -8183;
sin_rom[1453] = -8184;
sin_rom[1454] = -8185;
sin_rom[1455] = -8186;
sin_rom[1456] = -8187;
sin_rom[1457] = -8188;
sin_rom[1458] = -8189;
sin_rom[1459] = -8189;
sin_rom[1460] = -8190;
sin_rom[1461] = -8190;
sin_rom[1462] = -8191;
sin_rom[1463] = -8191;
sin_rom[1464] = -8191;
sin_rom[1465] = -8191;
sin_rom[1466] = -8191;
sin_rom[1467] = -8191;
sin_rom[1468] = -8191;
sin_rom[1469] = -8191;
sin_rom[1470] = -8191;
sin_rom[1471] = -8191;
sin_rom[1472] = -8190;
sin_rom[1473] = -8190;
sin_rom[1474] = -8189;
sin_rom[1475] = -8188;
sin_rom[1476] = -8187;
sin_rom[1477] = -8187;
sin_rom[1478] = -8186;
sin_rom[1479] = -8185;
sin_rom[1480] = -8183;
sin_rom[1481] = -8182;
sin_rom[1482] = -8181;
sin_rom[1483] = -8180;
sin_rom[1484] = -8178;
sin_rom[1485] = -8177;
sin_rom[1486] = -8175;
sin_rom[1487] = -8173;
sin_rom[1488] = -8171;
sin_rom[1489] = -8170;
sin_rom[1490] = -8168;
sin_rom[1491] = -8166;
sin_rom[1492] = -8163;
sin_rom[1493] = -8161;
sin_rom[1494] = -8159;
sin_rom[1495] = -8157;
sin_rom[1496] = -8154;
sin_rom[1497] = -8152;
sin_rom[1498] = -8149;
sin_rom[1499] = -8146;
sin_rom[1500] = -8143;
sin_rom[1501] = -8140;
sin_rom[1502] = -8137;
sin_rom[1503] = -8134;
sin_rom[1504] = -8131;
sin_rom[1505] = -8128;
sin_rom[1506] = -8125;
sin_rom[1507] = -8121;
sin_rom[1508] = -8118;
sin_rom[1509] = -8114;
sin_rom[1510] = -8111;
sin_rom[1511] = -8107;
sin_rom[1512] = -8103;
sin_rom[1513] = -8099;
sin_rom[1514] = -8095;
sin_rom[1515] = -8091;
sin_rom[1516] = -8087;
sin_rom[1517] = -8083;
sin_rom[1518] = -8078;
sin_rom[1519] = -8074;
sin_rom[1520] = -8070;
sin_rom[1521] = -8065;
sin_rom[1522] = -8060;
sin_rom[1523] = -8056;
sin_rom[1524] = -8051;
sin_rom[1525] = -8046;
sin_rom[1526] = -8041;
sin_rom[1527] = -8036;
sin_rom[1528] = -8031;
sin_rom[1529] = -8025;
sin_rom[1530] = -8020;
sin_rom[1531] = -8015;
sin_rom[1532] = -8009;
sin_rom[1533] = -8004;
sin_rom[1534] = -7998;
sin_rom[1535] = -7992;
sin_rom[1536] = -7986;
sin_rom[1537] = -7981;
sin_rom[1538] = -7975;
sin_rom[1539] = -7969;
sin_rom[1540] = -7962;
sin_rom[1541] = -7956;
sin_rom[1542] = -7950;
sin_rom[1543] = -7943;
sin_rom[1544] = -7937;
sin_rom[1545] = -7930;
sin_rom[1546] = -7924;
sin_rom[1547] = -7917;
sin_rom[1548] = -7910;
sin_rom[1549] = -7903;
sin_rom[1550] = -7896;
sin_rom[1551] = -7889;
sin_rom[1552] = -7882;
sin_rom[1553] = -7875;
sin_rom[1554] = -7868;
sin_rom[1555] = -7860;
sin_rom[1556] = -7853;
sin_rom[1557] = -7845;
sin_rom[1558] = -7838;
sin_rom[1559] = -7830;
sin_rom[1560] = -7822;
sin_rom[1561] = -7815;
sin_rom[1562] = -7807;
sin_rom[1563] = -7799;
sin_rom[1564] = -7790;
sin_rom[1565] = -7782;
sin_rom[1566] = -7774;
sin_rom[1567] = -7766;
sin_rom[1568] = -7757;
sin_rom[1569] = -7749;
sin_rom[1570] = -7740;
sin_rom[1571] = -7732;
sin_rom[1572] = -7723;
sin_rom[1573] = -7714;
sin_rom[1574] = -7705;
sin_rom[1575] = -7696;
sin_rom[1576] = -7687;
sin_rom[1577] = -7678;
sin_rom[1578] = -7669;
sin_rom[1579] = -7659;
sin_rom[1580] = -7650;
sin_rom[1581] = -7641;
sin_rom[1582] = -7631;
sin_rom[1583] = -7621;
sin_rom[1584] = -7612;
sin_rom[1585] = -7602;
sin_rom[1586] = -7592;
sin_rom[1587] = -7582;
sin_rom[1588] = -7572;
sin_rom[1589] = -7562;
sin_rom[1590] = -7552;
sin_rom[1591] = -7542;
sin_rom[1592] = -7531;
sin_rom[1593] = -7521;
sin_rom[1594] = -7511;
sin_rom[1595] = -7500;
sin_rom[1596] = -7489;
sin_rom[1597] = -7479;
sin_rom[1598] = -7468;
sin_rom[1599] = -7457;
sin_rom[1600] = -7446;
sin_rom[1601] = -7435;
sin_rom[1602] = -7424;
sin_rom[1603] = -7413;
sin_rom[1604] = -7402;
sin_rom[1605] = -7390;
sin_rom[1606] = -7379;
sin_rom[1607] = -7367;
sin_rom[1608] = -7356;
sin_rom[1609] = -7344;
sin_rom[1610] = -7333;
sin_rom[1611] = -7321;
sin_rom[1612] = -7309;
sin_rom[1613] = -7297;
sin_rom[1614] = -7285;
sin_rom[1615] = -7273;
sin_rom[1616] = -7261;
sin_rom[1617] = -7249;
sin_rom[1618] = -7236;
sin_rom[1619] = -7224;
sin_rom[1620] = -7211;
sin_rom[1621] = -7199;
sin_rom[1622] = -7186;
sin_rom[1623] = -7174;
sin_rom[1624] = -7161;
sin_rom[1625] = -7148;
sin_rom[1626] = -7135;
sin_rom[1627] = -7122;
sin_rom[1628] = -7109;
sin_rom[1629] = -7096;
sin_rom[1630] = -7083;
sin_rom[1631] = -7070;
sin_rom[1632] = -7056;
sin_rom[1633] = -7043;
sin_rom[1634] = -7029;
sin_rom[1635] = -7016;
sin_rom[1636] = -7002;
sin_rom[1637] = -6989;
sin_rom[1638] = -6975;
sin_rom[1639] = -6961;
sin_rom[1640] = -6947;
sin_rom[1641] = -6933;
sin_rom[1642] = -6919;
sin_rom[1643] = -6905;
sin_rom[1644] = -6891;
sin_rom[1645] = -6876;
sin_rom[1646] = -6862;
sin_rom[1647] = -6848;
sin_rom[1648] = -6833;
sin_rom[1649] = -6819;
sin_rom[1650] = -6804;
sin_rom[1651] = -6789;
sin_rom[1652] = -6774;
sin_rom[1653] = -6760;
sin_rom[1654] = -6745;
sin_rom[1655] = -6730;
sin_rom[1656] = -6715;
sin_rom[1657] = -6700;
sin_rom[1658] = -6684;
sin_rom[1659] = -6669;
sin_rom[1660] = -6654;
sin_rom[1661] = -6638;
sin_rom[1662] = -6623;
sin_rom[1663] = -6607;
sin_rom[1664] = -6592;
sin_rom[1665] = -6576;
sin_rom[1666] = -6560;
sin_rom[1667] = -6545;
sin_rom[1668] = -6529;
sin_rom[1669] = -6513;
sin_rom[1670] = -6497;
sin_rom[1671] = -6481;
sin_rom[1672] = -6465;
sin_rom[1673] = -6448;
sin_rom[1674] = -6432;
sin_rom[1675] = -6416;
sin_rom[1676] = -6399;
sin_rom[1677] = -6383;
sin_rom[1678] = -6366;
sin_rom[1679] = -6350;
sin_rom[1680] = -6333;
sin_rom[1681] = -6316;
sin_rom[1682] = -6300;
sin_rom[1683] = -6283;
sin_rom[1684] = -6266;
sin_rom[1685] = -6249;
sin_rom[1686] = -6232;
sin_rom[1687] = -6215;
sin_rom[1688] = -6198;
sin_rom[1689] = -6180;
sin_rom[1690] = -6163;
sin_rom[1691] = -6146;
sin_rom[1692] = -6128;
sin_rom[1693] = -6111;
sin_rom[1694] = -6093;
sin_rom[1695] = -6075;
sin_rom[1696] = -6058;
sin_rom[1697] = -6040;
sin_rom[1698] = -6022;
sin_rom[1699] = -6004;
sin_rom[1700] = -5986;
sin_rom[1701] = -5968;
sin_rom[1702] = -5950;
sin_rom[1703] = -5932;
sin_rom[1704] = -5914;
sin_rom[1705] = -5896;
sin_rom[1706] = -5877;
sin_rom[1707] = -5859;
sin_rom[1708] = -5841;
sin_rom[1709] = -5822;
sin_rom[1710] = -5804;
sin_rom[1711] = -5785;
sin_rom[1712] = -5766;
sin_rom[1713] = -5748;
sin_rom[1714] = -5729;
sin_rom[1715] = -5710;
sin_rom[1716] = -5691;
sin_rom[1717] = -5672;
sin_rom[1718] = -5653;
sin_rom[1719] = -5634;
sin_rom[1720] = -5615;
sin_rom[1721] = -5596;
sin_rom[1722] = -5576;
sin_rom[1723] = -5557;
sin_rom[1724] = -5538;
sin_rom[1725] = -5518;
sin_rom[1726] = -5499;
sin_rom[1727] = -5479;
sin_rom[1728] = -5460;
sin_rom[1729] = -5440;
sin_rom[1730] = -5420;
sin_rom[1731] = -5400;
sin_rom[1732] = -5381;
sin_rom[1733] = -5361;
sin_rom[1734] = -5341;
sin_rom[1735] = -5321;
sin_rom[1736] = -5301;
sin_rom[1737] = -5281;
sin_rom[1738] = -5261;
sin_rom[1739] = -5240;
sin_rom[1740] = -5220;
sin_rom[1741] = -5200;
sin_rom[1742] = -5179;
sin_rom[1743] = -5159;
sin_rom[1744] = -5139;
sin_rom[1745] = -5118;
sin_rom[1746] = -5097;
sin_rom[1747] = -5077;
sin_rom[1748] = -5056;
sin_rom[1749] = -5035;
sin_rom[1750] = -5015;
sin_rom[1751] = -4994;
sin_rom[1752] = -4973;
sin_rom[1753] = -4952;
sin_rom[1754] = -4931;
sin_rom[1755] = -4910;
sin_rom[1756] = -4889;
sin_rom[1757] = -4868;
sin_rom[1758] = -4846;
sin_rom[1759] = -4825;
sin_rom[1760] = -4804;
sin_rom[1761] = -4782;
sin_rom[1762] = -4761;
sin_rom[1763] = -4740;
sin_rom[1764] = -4718;
sin_rom[1765] = -4697;
sin_rom[1766] = -4675;
sin_rom[1767] = -4653;
sin_rom[1768] = -4632;
sin_rom[1769] = -4610;
sin_rom[1770] = -4588;
sin_rom[1771] = -4566;
sin_rom[1772] = -4544;
sin_rom[1773] = -4522;
sin_rom[1774] = -4500;
sin_rom[1775] = -4478;
sin_rom[1776] = -4456;
sin_rom[1777] = -4434;
sin_rom[1778] = -4412;
sin_rom[1779] = -4390;
sin_rom[1780] = -4368;
sin_rom[1781] = -4345;
sin_rom[1782] = -4323;
sin_rom[1783] = -4301;
sin_rom[1784] = -4278;
sin_rom[1785] = -4256;
sin_rom[1786] = -4233;
sin_rom[1787] = -4211;
sin_rom[1788] = -4188;
sin_rom[1789] = -4165;
sin_rom[1790] = -4143;
sin_rom[1791] = -4120;
sin_rom[1792] = -4097;
sin_rom[1793] = -4074;
sin_rom[1794] = -4052;
sin_rom[1795] = -4029;
sin_rom[1796] = -4006;
sin_rom[1797] = -3983;
sin_rom[1798] = -3960;
sin_rom[1799] = -3937;
sin_rom[1800] = -3913;
sin_rom[1801] = -3890;
sin_rom[1802] = -3867;
sin_rom[1803] = -3844;
sin_rom[1804] = -3821;
sin_rom[1805] = -3797;
sin_rom[1806] = -3774;
sin_rom[1807] = -3751;
sin_rom[1808] = -3727;
sin_rom[1809] = -3704;
sin_rom[1810] = -3680;
sin_rom[1811] = -3657;
sin_rom[1812] = -3633;
sin_rom[1813] = -3609;
sin_rom[1814] = -3586;
sin_rom[1815] = -3562;
sin_rom[1816] = -3538;
sin_rom[1817] = -3515;
sin_rom[1818] = -3491;
sin_rom[1819] = -3467;
sin_rom[1820] = -3443;
sin_rom[1821] = -3419;
sin_rom[1822] = -3395;
sin_rom[1823] = -3371;
sin_rom[1824] = -3347;
sin_rom[1825] = -3323;
sin_rom[1826] = -3299;
sin_rom[1827] = -3275;
sin_rom[1828] = -3251;
sin_rom[1829] = -3227;
sin_rom[1830] = -3203;
sin_rom[1831] = -3178;
sin_rom[1832] = -3154;
sin_rom[1833] = -3130;
sin_rom[1834] = -3105;
sin_rom[1835] = -3081;
sin_rom[1836] = -3057;
sin_rom[1837] = -3032;
sin_rom[1838] = -3008;
sin_rom[1839] = -2983;
sin_rom[1840] = -2959;
sin_rom[1841] = -2934;
sin_rom[1842] = -2909;
sin_rom[1843] = -2885;
sin_rom[1844] = -2860;
sin_rom[1845] = -2835;
sin_rom[1846] = -2811;
sin_rom[1847] = -2786;
sin_rom[1848] = -2761;
sin_rom[1849] = -2736;
sin_rom[1850] = -2712;
sin_rom[1851] = -2687;
sin_rom[1852] = -2662;
sin_rom[1853] = -2637;
sin_rom[1854] = -2612;
sin_rom[1855] = -2587;
sin_rom[1856] = -2562;
sin_rom[1857] = -2537;
sin_rom[1858] = -2512;
sin_rom[1859] = -2487;
sin_rom[1860] = -2462;
sin_rom[1861] = -2437;
sin_rom[1862] = -2412;
sin_rom[1863] = -2386;
sin_rom[1864] = -2361;
sin_rom[1865] = -2336;
sin_rom[1866] = -2311;
sin_rom[1867] = -2285;
sin_rom[1868] = -2260;
sin_rom[1869] = -2235;
sin_rom[1870] = -2209;
sin_rom[1871] = -2184;
sin_rom[1872] = -2159;
sin_rom[1873] = -2133;
sin_rom[1874] = -2108;
sin_rom[1875] = -2082;
sin_rom[1876] = -2057;
sin_rom[1877] = -2031;
sin_rom[1878] = -2006;
sin_rom[1879] = -1980;
sin_rom[1880] = -1955;
sin_rom[1881] = -1929;
sin_rom[1882] = -1904;
sin_rom[1883] = -1878;
sin_rom[1884] = -1852;
sin_rom[1885] = -1827;
sin_rom[1886] = -1801;
sin_rom[1887] = -1775;
sin_rom[1888] = -1750;
sin_rom[1889] = -1724;
sin_rom[1890] = -1698;
sin_rom[1891] = -1672;
sin_rom[1892] = -1647;
sin_rom[1893] = -1621;
sin_rom[1894] = -1595;
sin_rom[1895] = -1569;
sin_rom[1896] = -1543;
sin_rom[1897] = -1517;
sin_rom[1898] = -1492;
sin_rom[1899] = -1466;
sin_rom[1900] = -1440;
sin_rom[1901] = -1414;
sin_rom[1902] = -1388;
sin_rom[1903] = -1362;
sin_rom[1904] = -1336;
sin_rom[1905] = -1310;
sin_rom[1906] = -1284;
sin_rom[1907] = -1258;
sin_rom[1908] = -1232;
sin_rom[1909] = -1206;
sin_rom[1910] = -1180;
sin_rom[1911] = -1154;
sin_rom[1912] = -1128;
sin_rom[1913] = -1102;
sin_rom[1914] = -1076;
sin_rom[1915] = -1050;
sin_rom[1916] = -1023;
sin_rom[1917] = -997;
sin_rom[1918] = -971;
sin_rom[1919] = -945;
sin_rom[1920] = -919;
sin_rom[1921] = -893;
sin_rom[1922] = -866;
sin_rom[1923] = -840;
sin_rom[1924] = -814;
sin_rom[1925] = -788;
sin_rom[1926] = -762;
sin_rom[1927] = -735;
sin_rom[1928] = -709;
sin_rom[1929] = -683;
sin_rom[1930] = -657;
sin_rom[1931] = -631;
sin_rom[1932] = -604;
sin_rom[1933] = -578;
sin_rom[1934] = -552;
sin_rom[1935] = -525;
sin_rom[1936] = -499;
sin_rom[1937] = -473;
sin_rom[1938] = -447;
sin_rom[1939] = -420;
sin_rom[1940] = -394;
sin_rom[1941] = -368;
sin_rom[1942] = -341;
sin_rom[1943] = -315;
sin_rom[1944] = -289;
sin_rom[1945] = -263;
sin_rom[1946] = -236;
sin_rom[1947] = -210;
sin_rom[1948] = -184;
sin_rom[1949] = -157;
sin_rom[1950] = -131;
sin_rom[1951] = -105;
sin_rom[1952] = -78;
sin_rom[1953] = -52;
end


reg [18:0]addr = phase*500000/360;

always@(posedge clk)begin
    if(addr+freq<500000)
        addr<=addr+freq;
    else
        addr<=addr+freq-500000;
    dds_o<=sin_rom[addr[18:8]];
end

endmodule

module dds_p(
input clk,
input [13:0]freq,
input [13:0]phase,
output reg signed [13:0]dds_o 
);


reg signed [13:0] sin_rom [0:1953];
initial begin
sin_rom[0] = 0;
sin_rom[1] = 26;
sin_rom[2] = 52;
sin_rom[3] = 78;
sin_rom[4] = 105;
sin_rom[5] = 131;
sin_rom[6] = 157;
sin_rom[7] = 184;
sin_rom[8] = 210;
sin_rom[9] = 236;
sin_rom[10] = 263;
sin_rom[11] = 289;
sin_rom[12] = 315;
sin_rom[13] = 342;
sin_rom[14] = 368;
sin_rom[15] = 394;
sin_rom[16] = 421;
sin_rom[17] = 447;
sin_rom[18] = 473;
sin_rom[19] = 499;
sin_rom[20] = 526;
sin_rom[21] = 552;
sin_rom[22] = 578;
sin_rom[23] = 605;
sin_rom[24] = 631;
sin_rom[25] = 657;
sin_rom[26] = 683;
sin_rom[27] = 709;
sin_rom[28] = 736;
sin_rom[29] = 762;
sin_rom[30] = 788;
sin_rom[31] = 814;
sin_rom[32] = 841;
sin_rom[33] = 867;
sin_rom[34] = 893;
sin_rom[35] = 919;
sin_rom[36] = 945;
sin_rom[37] = 971;
sin_rom[38] = 997;
sin_rom[39] = 1024;
sin_rom[40] = 1050;
sin_rom[41] = 1076;
sin_rom[42] = 1102;
sin_rom[43] = 1128;
sin_rom[44] = 1154;
sin_rom[45] = 1180;
sin_rom[46] = 1206;
sin_rom[47] = 1232;
sin_rom[48] = 1258;
sin_rom[49] = 1284;
sin_rom[50] = 1310;
sin_rom[51] = 1336;
sin_rom[52] = 1362;
sin_rom[53] = 1388;
sin_rom[54] = 1414;
sin_rom[55] = 1440;
sin_rom[56] = 1466;
sin_rom[57] = 1492;
sin_rom[58] = 1518;
sin_rom[59] = 1544;
sin_rom[60] = 1569;
sin_rom[61] = 1595;
sin_rom[62] = 1621;
sin_rom[63] = 1647;
sin_rom[64] = 1673;
sin_rom[65] = 1698;
sin_rom[66] = 1724;
sin_rom[67] = 1750;
sin_rom[68] = 1776;
sin_rom[69] = 1801;
sin_rom[70] = 1827;
sin_rom[71] = 1853;
sin_rom[72] = 1878;
sin_rom[73] = 1904;
sin_rom[74] = 1929;
sin_rom[75] = 1955;
sin_rom[76] = 1981;
sin_rom[77] = 2006;
sin_rom[78] = 2032;
sin_rom[79] = 2057;
sin_rom[80] = 2083;
sin_rom[81] = 2108;
sin_rom[82] = 2134;
sin_rom[83] = 2159;
sin_rom[84] = 2184;
sin_rom[85] = 2210;
sin_rom[86] = 2235;
sin_rom[87] = 2260;
sin_rom[88] = 2286;
sin_rom[89] = 2311;
sin_rom[90] = 2336;
sin_rom[91] = 2361;
sin_rom[92] = 2387;
sin_rom[93] = 2412;
sin_rom[94] = 2437;
sin_rom[95] = 2462;
sin_rom[96] = 2487;
sin_rom[97] = 2512;
sin_rom[98] = 2537;
sin_rom[99] = 2562;
sin_rom[100] = 2587;
sin_rom[101] = 2612;
sin_rom[102] = 2637;
sin_rom[103] = 2662;
sin_rom[104] = 2687;
sin_rom[105] = 2712;
sin_rom[106] = 2737;
sin_rom[107] = 2761;
sin_rom[108] = 2786;
sin_rom[109] = 2811;
sin_rom[110] = 2836;
sin_rom[111] = 2860;
sin_rom[112] = 2885;
sin_rom[113] = 2910;
sin_rom[114] = 2934;
sin_rom[115] = 2959;
sin_rom[116] = 2983;
sin_rom[117] = 3008;
sin_rom[118] = 3032;
sin_rom[119] = 3057;
sin_rom[120] = 3081;
sin_rom[121] = 3106;
sin_rom[122] = 3130;
sin_rom[123] = 3154;
sin_rom[124] = 3178;
sin_rom[125] = 3203;
sin_rom[126] = 3227;
sin_rom[127] = 3251;
sin_rom[128] = 3275;
sin_rom[129] = 3299;
sin_rom[130] = 3323;
sin_rom[131] = 3348;
sin_rom[132] = 3372;
sin_rom[133] = 3396;
sin_rom[134] = 3419;
sin_rom[135] = 3443;
sin_rom[136] = 3467;
sin_rom[137] = 3491;
sin_rom[138] = 3515;
sin_rom[139] = 3539;
sin_rom[140] = 3562;
sin_rom[141] = 3586;
sin_rom[142] = 3610;
sin_rom[143] = 3633;
sin_rom[144] = 3657;
sin_rom[145] = 3680;
sin_rom[146] = 3704;
sin_rom[147] = 3727;
sin_rom[148] = 3751;
sin_rom[149] = 3774;
sin_rom[150] = 3798;
sin_rom[151] = 3821;
sin_rom[152] = 3844;
sin_rom[153] = 3867;
sin_rom[154] = 3891;
sin_rom[155] = 3914;
sin_rom[156] = 3937;
sin_rom[157] = 3960;
sin_rom[158] = 3983;
sin_rom[159] = 4006;
sin_rom[160] = 4029;
sin_rom[161] = 4052;
sin_rom[162] = 4075;
sin_rom[163] = 4097;
sin_rom[164] = 4120;
sin_rom[165] = 4143;
sin_rom[166] = 4166;
sin_rom[167] = 4188;
sin_rom[168] = 4211;
sin_rom[169] = 4233;
sin_rom[170] = 4256;
sin_rom[171] = 4278;
sin_rom[172] = 4301;
sin_rom[173] = 4323;
sin_rom[174] = 4346;
sin_rom[175] = 4368;
sin_rom[176] = 4390;
sin_rom[177] = 4412;
sin_rom[178] = 4434;
sin_rom[179] = 4457;
sin_rom[180] = 4479;
sin_rom[181] = 4501;
sin_rom[182] = 4523;
sin_rom[183] = 4545;
sin_rom[184] = 4566;
sin_rom[185] = 4588;
sin_rom[186] = 4610;
sin_rom[187] = 4632;
sin_rom[188] = 4654;
sin_rom[189] = 4675;
sin_rom[190] = 4697;
sin_rom[191] = 4718;
sin_rom[192] = 4740;
sin_rom[193] = 4761;
sin_rom[194] = 4783;
sin_rom[195] = 4804;
sin_rom[196] = 4825;
sin_rom[197] = 4847;
sin_rom[198] = 4868;
sin_rom[199] = 4889;
sin_rom[200] = 4910;
sin_rom[201] = 4931;
sin_rom[202] = 4952;
sin_rom[203] = 4973;
sin_rom[204] = 4994;
sin_rom[205] = 5015;
sin_rom[206] = 5036;
sin_rom[207] = 5056;
sin_rom[208] = 5077;
sin_rom[209] = 5098;
sin_rom[210] = 5118;
sin_rom[211] = 5139;
sin_rom[212] = 5159;
sin_rom[213] = 5180;
sin_rom[214] = 5200;
sin_rom[215] = 5220;
sin_rom[216] = 5241;
sin_rom[217] = 5261;
sin_rom[218] = 5281;
sin_rom[219] = 5301;
sin_rom[220] = 5321;
sin_rom[221] = 5341;
sin_rom[222] = 5361;
sin_rom[223] = 5381;
sin_rom[224] = 5401;
sin_rom[225] = 5420;
sin_rom[226] = 5440;
sin_rom[227] = 5460;
sin_rom[228] = 5479;
sin_rom[229] = 5499;
sin_rom[230] = 5518;
sin_rom[231] = 5538;
sin_rom[232] = 5557;
sin_rom[233] = 5577;
sin_rom[234] = 5596;
sin_rom[235] = 5615;
sin_rom[236] = 5634;
sin_rom[237] = 5653;
sin_rom[238] = 5672;
sin_rom[239] = 5691;
sin_rom[240] = 5710;
sin_rom[241] = 5729;
sin_rom[242] = 5748;
sin_rom[243] = 5766;
sin_rom[244] = 5785;
sin_rom[245] = 5804;
sin_rom[246] = 5822;
sin_rom[247] = 5841;
sin_rom[248] = 5859;
sin_rom[249] = 5878;
sin_rom[250] = 5896;
sin_rom[251] = 5914;
sin_rom[252] = 5932;
sin_rom[253] = 5950;
sin_rom[254] = 5969;
sin_rom[255] = 5987;
sin_rom[256] = 6004;
sin_rom[257] = 6022;
sin_rom[258] = 6040;
sin_rom[259] = 6058;
sin_rom[260] = 6076;
sin_rom[261] = 6093;
sin_rom[262] = 6111;
sin_rom[263] = 6128;
sin_rom[264] = 6146;
sin_rom[265] = 6163;
sin_rom[266] = 6180;
sin_rom[267] = 6198;
sin_rom[268] = 6215;
sin_rom[269] = 6232;
sin_rom[270] = 6249;
sin_rom[271] = 6266;
sin_rom[272] = 6283;
sin_rom[273] = 6300;
sin_rom[274] = 6317;
sin_rom[275] = 6333;
sin_rom[276] = 6350;
sin_rom[277] = 6367;
sin_rom[278] = 6383;
sin_rom[279] = 6400;
sin_rom[280] = 6416;
sin_rom[281] = 6432;
sin_rom[282] = 6449;
sin_rom[283] = 6465;
sin_rom[284] = 6481;
sin_rom[285] = 6497;
sin_rom[286] = 6513;
sin_rom[287] = 6529;
sin_rom[288] = 6545;
sin_rom[289] = 6561;
sin_rom[290] = 6576;
sin_rom[291] = 6592;
sin_rom[292] = 6608;
sin_rom[293] = 6623;
sin_rom[294] = 6639;
sin_rom[295] = 6654;
sin_rom[296] = 6669;
sin_rom[297] = 6685;
sin_rom[298] = 6700;
sin_rom[299] = 6715;
sin_rom[300] = 6730;
sin_rom[301] = 6745;
sin_rom[302] = 6760;
sin_rom[303] = 6775;
sin_rom[304] = 6789;
sin_rom[305] = 6804;
sin_rom[306] = 6819;
sin_rom[307] = 6833;
sin_rom[308] = 6848;
sin_rom[309] = 6862;
sin_rom[310] = 6876;
sin_rom[311] = 6891;
sin_rom[312] = 6905;
sin_rom[313] = 6919;
sin_rom[314] = 6933;
sin_rom[315] = 6947;
sin_rom[316] = 6961;
sin_rom[317] = 6975;
sin_rom[318] = 6989;
sin_rom[319] = 7002;
sin_rom[320] = 7016;
sin_rom[321] = 7030;
sin_rom[322] = 7043;
sin_rom[323] = 7056;
sin_rom[324] = 7070;
sin_rom[325] = 7083;
sin_rom[326] = 7096;
sin_rom[327] = 7109;
sin_rom[328] = 7122;
sin_rom[329] = 7135;
sin_rom[330] = 7148;
sin_rom[331] = 7161;
sin_rom[332] = 7174;
sin_rom[333] = 7186;
sin_rom[334] = 7199;
sin_rom[335] = 7212;
sin_rom[336] = 7224;
sin_rom[337] = 7236;
sin_rom[338] = 7249;
sin_rom[339] = 7261;
sin_rom[340] = 7273;
sin_rom[341] = 7285;
sin_rom[342] = 7297;
sin_rom[343] = 7309;
sin_rom[344] = 7321;
sin_rom[345] = 7333;
sin_rom[346] = 7344;
sin_rom[347] = 7356;
sin_rom[348] = 7368;
sin_rom[349] = 7379;
sin_rom[350] = 7390;
sin_rom[351] = 7402;
sin_rom[352] = 7413;
sin_rom[353] = 7424;
sin_rom[354] = 7435;
sin_rom[355] = 7446;
sin_rom[356] = 7457;
sin_rom[357] = 7468;
sin_rom[358] = 7479;
sin_rom[359] = 7490;
sin_rom[360] = 7500;
sin_rom[361] = 7511;
sin_rom[362] = 7521;
sin_rom[363] = 7532;
sin_rom[364] = 7542;
sin_rom[365] = 7552;
sin_rom[366] = 7562;
sin_rom[367] = 7572;
sin_rom[368] = 7582;
sin_rom[369] = 7592;
sin_rom[370] = 7602;
sin_rom[371] = 7612;
sin_rom[372] = 7622;
sin_rom[373] = 7631;
sin_rom[374] = 7641;
sin_rom[375] = 7650;
sin_rom[376] = 7660;
sin_rom[377] = 7669;
sin_rom[378] = 7678;
sin_rom[379] = 7687;
sin_rom[380] = 7696;
sin_rom[381] = 7705;
sin_rom[382] = 7714;
sin_rom[383] = 7723;
sin_rom[384] = 7732;
sin_rom[385] = 7740;
sin_rom[386] = 7749;
sin_rom[387] = 7757;
sin_rom[388] = 7766;
sin_rom[389] = 7774;
sin_rom[390] = 7782;
sin_rom[391] = 7791;
sin_rom[392] = 7799;
sin_rom[393] = 7807;
sin_rom[394] = 7815;
sin_rom[395] = 7822;
sin_rom[396] = 7830;
sin_rom[397] = 7838;
sin_rom[398] = 7846;
sin_rom[399] = 7853;
sin_rom[400] = 7861;
sin_rom[401] = 7868;
sin_rom[402] = 7875;
sin_rom[403] = 7882;
sin_rom[404] = 7890;
sin_rom[405] = 7897;
sin_rom[406] = 7904;
sin_rom[407] = 7910;
sin_rom[408] = 7917;
sin_rom[409] = 7924;
sin_rom[410] = 7931;
sin_rom[411] = 7937;
sin_rom[412] = 7944;
sin_rom[413] = 7950;
sin_rom[414] = 7956;
sin_rom[415] = 7962;
sin_rom[416] = 7969;
sin_rom[417] = 7975;
sin_rom[418] = 7981;
sin_rom[419] = 7987;
sin_rom[420] = 7992;
sin_rom[421] = 7998;
sin_rom[422] = 8004;
sin_rom[423] = 8009;
sin_rom[424] = 8015;
sin_rom[425] = 8020;
sin_rom[426] = 8025;
sin_rom[427] = 8031;
sin_rom[428] = 8036;
sin_rom[429] = 8041;
sin_rom[430] = 8046;
sin_rom[431] = 8051;
sin_rom[432] = 8056;
sin_rom[433] = 8060;
sin_rom[434] = 8065;
sin_rom[435] = 8070;
sin_rom[436] = 8074;
sin_rom[437] = 8078;
sin_rom[438] = 8083;
sin_rom[439] = 8087;
sin_rom[440] = 8091;
sin_rom[441] = 8095;
sin_rom[442] = 8099;
sin_rom[443] = 8103;
sin_rom[444] = 8107;
sin_rom[445] = 8111;
sin_rom[446] = 8114;
sin_rom[447] = 8118;
sin_rom[448] = 8121;
sin_rom[449] = 8125;
sin_rom[450] = 8128;
sin_rom[451] = 8131;
sin_rom[452] = 8134;
sin_rom[453] = 8137;
sin_rom[454] = 8140;
sin_rom[455] = 8143;
sin_rom[456] = 8146;
sin_rom[457] = 8149;
sin_rom[458] = 8152;
sin_rom[459] = 8154;
sin_rom[460] = 8157;
sin_rom[461] = 8159;
sin_rom[462] = 8161;
sin_rom[463] = 8163;
sin_rom[464] = 8166;
sin_rom[465] = 8168;
sin_rom[466] = 8170;
sin_rom[467] = 8171;
sin_rom[468] = 8173;
sin_rom[469] = 8175;
sin_rom[470] = 8177;
sin_rom[471] = 8178;
sin_rom[472] = 8180;
sin_rom[473] = 8181;
sin_rom[474] = 8182;
sin_rom[475] = 8184;
sin_rom[476] = 8185;
sin_rom[477] = 8186;
sin_rom[478] = 8187;
sin_rom[479] = 8187;
sin_rom[480] = 8188;
sin_rom[481] = 8189;
sin_rom[482] = 8190;
sin_rom[483] = 8190;
sin_rom[484] = 8191;
sin_rom[485] = 8191;
sin_rom[486] = 8191;
sin_rom[487] = 8191;
sin_rom[488] = 8191;
sin_rom[489] = 8191;
sin_rom[490] = 8191;
sin_rom[491] = 8191;
sin_rom[492] = 8191;
sin_rom[493] = 8191;
sin_rom[494] = 8190;
sin_rom[495] = 8190;
sin_rom[496] = 8189;
sin_rom[497] = 8189;
sin_rom[498] = 8188;
sin_rom[499] = 8187;
sin_rom[500] = 8186;
sin_rom[501] = 8185;
sin_rom[502] = 8184;
sin_rom[503] = 8183;
sin_rom[504] = 8182;
sin_rom[505] = 8180;
sin_rom[506] = 8179;
sin_rom[507] = 8177;
sin_rom[508] = 8176;
sin_rom[509] = 8174;
sin_rom[510] = 8172;
sin_rom[511] = 8171;
sin_rom[512] = 8169;
sin_rom[513] = 8167;
sin_rom[514] = 8165;
sin_rom[515] = 8162;
sin_rom[516] = 8160;
sin_rom[517] = 8158;
sin_rom[518] = 8155;
sin_rom[519] = 8153;
sin_rom[520] = 8150;
sin_rom[521] = 8148;
sin_rom[522] = 8145;
sin_rom[523] = 8142;
sin_rom[524] = 8139;
sin_rom[525] = 8136;
sin_rom[526] = 8133;
sin_rom[527] = 8130;
sin_rom[528] = 8126;
sin_rom[529] = 8123;
sin_rom[530] = 8120;
sin_rom[531] = 8116;
sin_rom[532] = 8112;
sin_rom[533] = 8109;
sin_rom[534] = 8105;
sin_rom[535] = 8101;
sin_rom[536] = 8097;
sin_rom[537] = 8093;
sin_rom[538] = 8089;
sin_rom[539] = 8085;
sin_rom[540] = 8081;
sin_rom[541] = 8076;
sin_rom[542] = 8072;
sin_rom[543] = 8067;
sin_rom[544] = 8063;
sin_rom[545] = 8058;
sin_rom[546] = 8053;
sin_rom[547] = 8048;
sin_rom[548] = 8043;
sin_rom[549] = 8038;
sin_rom[550] = 8033;
sin_rom[551] = 8028;
sin_rom[552] = 8023;
sin_rom[553] = 8017;
sin_rom[554] = 8012;
sin_rom[555] = 8006;
sin_rom[556] = 8001;
sin_rom[557] = 7995;
sin_rom[558] = 7989;
sin_rom[559] = 7984;
sin_rom[560] = 7978;
sin_rom[561] = 7972;
sin_rom[562] = 7966;
sin_rom[563] = 7959;
sin_rom[564] = 7953;
sin_rom[565] = 7947;
sin_rom[566] = 7940;
sin_rom[567] = 7934;
sin_rom[568] = 7927;
sin_rom[569] = 7921;
sin_rom[570] = 7914;
sin_rom[571] = 7907;
sin_rom[572] = 7900;
sin_rom[573] = 7893;
sin_rom[574] = 7886;
sin_rom[575] = 7879;
sin_rom[576] = 7872;
sin_rom[577] = 7864;
sin_rom[578] = 7857;
sin_rom[579] = 7849;
sin_rom[580] = 7842;
sin_rom[581] = 7834;
sin_rom[582] = 7826;
sin_rom[583] = 7819;
sin_rom[584] = 7811;
sin_rom[585] = 7803;
sin_rom[586] = 7795;
sin_rom[587] = 7786;
sin_rom[588] = 7778;
sin_rom[589] = 7770;
sin_rom[590] = 7762;
sin_rom[591] = 7753;
sin_rom[592] = 7745;
sin_rom[593] = 7736;
sin_rom[594] = 7727;
sin_rom[595] = 7718;
sin_rom[596] = 7710;
sin_rom[597] = 7701;
sin_rom[598] = 7692;
sin_rom[599] = 7683;
sin_rom[600] = 7673;
sin_rom[601] = 7664;
sin_rom[602] = 7655;
sin_rom[603] = 7645;
sin_rom[604] = 7636;
sin_rom[605] = 7626;
sin_rom[606] = 7617;
sin_rom[607] = 7607;
sin_rom[608] = 7597;
sin_rom[609] = 7587;
sin_rom[610] = 7577;
sin_rom[611] = 7567;
sin_rom[612] = 7557;
sin_rom[613] = 7547;
sin_rom[614] = 7537;
sin_rom[615] = 7526;
sin_rom[616] = 7516;
sin_rom[617] = 7505;
sin_rom[618] = 7495;
sin_rom[619] = 7484;
sin_rom[620] = 7473;
sin_rom[621] = 7463;
sin_rom[622] = 7452;
sin_rom[623] = 7441;
sin_rom[624] = 7430;
sin_rom[625] = 7419;
sin_rom[626] = 7407;
sin_rom[627] = 7396;
sin_rom[628] = 7385;
sin_rom[629] = 7373;
sin_rom[630] = 7362;
sin_rom[631] = 7350;
sin_rom[632] = 7339;
sin_rom[633] = 7327;
sin_rom[634] = 7315;
sin_rom[635] = 7303;
sin_rom[636] = 7291;
sin_rom[637] = 7279;
sin_rom[638] = 7267;
sin_rom[639] = 7255;
sin_rom[640] = 7243;
sin_rom[641] = 7230;
sin_rom[642] = 7218;
sin_rom[643] = 7205;
sin_rom[644] = 7193;
sin_rom[645] = 7180;
sin_rom[646] = 7167;
sin_rom[647] = 7155;
sin_rom[648] = 7142;
sin_rom[649] = 7129;
sin_rom[650] = 7116;
sin_rom[651] = 7103;
sin_rom[652] = 7090;
sin_rom[653] = 7076;
sin_rom[654] = 7063;
sin_rom[655] = 7050;
sin_rom[656] = 7036;
sin_rom[657] = 7023;
sin_rom[658] = 7009;
sin_rom[659] = 6995;
sin_rom[660] = 6982;
sin_rom[661] = 6968;
sin_rom[662] = 6954;
sin_rom[663] = 6940;
sin_rom[664] = 6926;
sin_rom[665] = 6912;
sin_rom[666] = 6898;
sin_rom[667] = 6884;
sin_rom[668] = 6869;
sin_rom[669] = 6855;
sin_rom[670] = 6840;
sin_rom[671] = 6826;
sin_rom[672] = 6811;
sin_rom[673] = 6797;
sin_rom[674] = 6782;
sin_rom[675] = 6767;
sin_rom[676] = 6752;
sin_rom[677] = 6737;
sin_rom[678] = 6722;
sin_rom[679] = 6707;
sin_rom[680] = 6692;
sin_rom[681] = 6677;
sin_rom[682] = 6662;
sin_rom[683] = 6646;
sin_rom[684] = 6631;
sin_rom[685] = 6615;
sin_rom[686] = 6600;
sin_rom[687] = 6584;
sin_rom[688] = 6568;
sin_rom[689] = 6553;
sin_rom[690] = 6537;
sin_rom[691] = 6521;
sin_rom[692] = 6505;
sin_rom[693] = 6489;
sin_rom[694] = 6473;
sin_rom[695] = 6457;
sin_rom[696] = 6440;
sin_rom[697] = 6424;
sin_rom[698] = 6408;
sin_rom[699] = 6391;
sin_rom[700] = 6375;
sin_rom[701] = 6358;
sin_rom[702] = 6342;
sin_rom[703] = 6325;
sin_rom[704] = 6308;
sin_rom[705] = 6291;
sin_rom[706] = 6274;
sin_rom[707] = 6257;
sin_rom[708] = 6240;
sin_rom[709] = 6223;
sin_rom[710] = 6206;
sin_rom[711] = 6189;
sin_rom[712] = 6172;
sin_rom[713] = 6154;
sin_rom[714] = 6137;
sin_rom[715] = 6119;
sin_rom[716] = 6102;
sin_rom[717] = 6084;
sin_rom[718] = 6067;
sin_rom[719] = 6049;
sin_rom[720] = 6031;
sin_rom[721] = 6013;
sin_rom[722] = 5995;
sin_rom[723] = 5977;
sin_rom[724] = 5959;
sin_rom[725] = 5941;
sin_rom[726] = 5923;
sin_rom[727] = 5905;
sin_rom[728] = 5887;
sin_rom[729] = 5868;
sin_rom[730] = 5850;
sin_rom[731] = 5831;
sin_rom[732] = 5813;
sin_rom[733] = 5794;
sin_rom[734] = 5776;
sin_rom[735] = 5757;
sin_rom[736] = 5738;
sin_rom[737] = 5719;
sin_rom[738] = 5701;
sin_rom[739] = 5682;
sin_rom[740] = 5663;
sin_rom[741] = 5644;
sin_rom[742] = 5624;
sin_rom[743] = 5605;
sin_rom[744] = 5586;
sin_rom[745] = 5567;
sin_rom[746] = 5547;
sin_rom[747] = 5528;
sin_rom[748] = 5509;
sin_rom[749] = 5489;
sin_rom[750] = 5470;
sin_rom[751] = 5450;
sin_rom[752] = 5430;
sin_rom[753] = 5410;
sin_rom[754] = 5391;
sin_rom[755] = 5371;
sin_rom[756] = 5351;
sin_rom[757] = 5331;
sin_rom[758] = 5311;
sin_rom[759] = 5291;
sin_rom[760] = 5271;
sin_rom[761] = 5251;
sin_rom[762] = 5230;
sin_rom[763] = 5210;
sin_rom[764] = 5190;
sin_rom[765] = 5169;
sin_rom[766] = 5149;
sin_rom[767] = 5128;
sin_rom[768] = 5108;
sin_rom[769] = 5087;
sin_rom[770] = 5067;
sin_rom[771] = 5046;
sin_rom[772] = 5025;
sin_rom[773] = 5004;
sin_rom[774] = 4983;
sin_rom[775] = 4962;
sin_rom[776] = 4941;
sin_rom[777] = 4920;
sin_rom[778] = 4899;
sin_rom[779] = 4878;
sin_rom[780] = 4857;
sin_rom[781] = 4836;
sin_rom[782] = 4815;
sin_rom[783] = 4793;
sin_rom[784] = 4772;
sin_rom[785] = 4750;
sin_rom[786] = 4729;
sin_rom[787] = 4707;
sin_rom[788] = 4686;
sin_rom[789] = 4664;
sin_rom[790] = 4643;
sin_rom[791] = 4621;
sin_rom[792] = 4599;
sin_rom[793] = 4577;
sin_rom[794] = 4555;
sin_rom[795] = 4534;
sin_rom[796] = 4512;
sin_rom[797] = 4490;
sin_rom[798] = 4468;
sin_rom[799] = 4445;
sin_rom[800] = 4423;
sin_rom[801] = 4401;
sin_rom[802] = 4379;
sin_rom[803] = 4357;
sin_rom[804] = 4334;
sin_rom[805] = 4312;
sin_rom[806] = 4290;
sin_rom[807] = 4267;
sin_rom[808] = 4245;
sin_rom[809] = 4222;
sin_rom[810] = 4199;
sin_rom[811] = 4177;
sin_rom[812] = 4154;
sin_rom[813] = 4131;
sin_rom[814] = 4109;
sin_rom[815] = 4086;
sin_rom[816] = 4063;
sin_rom[817] = 4040;
sin_rom[818] = 4017;
sin_rom[819] = 3994;
sin_rom[820] = 3971;
sin_rom[821] = 3948;
sin_rom[822] = 3925;
sin_rom[823] = 3902;
sin_rom[824] = 3879;
sin_rom[825] = 3856;
sin_rom[826] = 3832;
sin_rom[827] = 3809;
sin_rom[828] = 3786;
sin_rom[829] = 3762;
sin_rom[830] = 3739;
sin_rom[831] = 3716;
sin_rom[832] = 3692;
sin_rom[833] = 3669;
sin_rom[834] = 3645;
sin_rom[835] = 3621;
sin_rom[836] = 3598;
sin_rom[837] = 3574;
sin_rom[838] = 3550;
sin_rom[839] = 3527;
sin_rom[840] = 3503;
sin_rom[841] = 3479;
sin_rom[842] = 3455;
sin_rom[843] = 3431;
sin_rom[844] = 3407;
sin_rom[845] = 3383;
sin_rom[846] = 3359;
sin_rom[847] = 3335;
sin_rom[848] = 3311;
sin_rom[849] = 3287;
sin_rom[850] = 3263;
sin_rom[851] = 3239;
sin_rom[852] = 3215;
sin_rom[853] = 3191;
sin_rom[854] = 3166;
sin_rom[855] = 3142;
sin_rom[856] = 3118;
sin_rom[857] = 3093;
sin_rom[858] = 3069;
sin_rom[859] = 3044;
sin_rom[860] = 3020;
sin_rom[861] = 2995;
sin_rom[862] = 2971;
sin_rom[863] = 2946;
sin_rom[864] = 2922;
sin_rom[865] = 2897;
sin_rom[866] = 2873;
sin_rom[867] = 2848;
sin_rom[868] = 2823;
sin_rom[869] = 2798;
sin_rom[870] = 2774;
sin_rom[871] = 2749;
sin_rom[872] = 2724;
sin_rom[873] = 2699;
sin_rom[874] = 2674;
sin_rom[875] = 2650;
sin_rom[876] = 2625;
sin_rom[877] = 2600;
sin_rom[878] = 2575;
sin_rom[879] = 2550;
sin_rom[880] = 2525;
sin_rom[881] = 2500;
sin_rom[882] = 2474;
sin_rom[883] = 2449;
sin_rom[884] = 2424;
sin_rom[885] = 2399;
sin_rom[886] = 2374;
sin_rom[887] = 2349;
sin_rom[888] = 2323;
sin_rom[889] = 2298;
sin_rom[890] = 2273;
sin_rom[891] = 2248;
sin_rom[892] = 2222;
sin_rom[893] = 2197;
sin_rom[894] = 2172;
sin_rom[895] = 2146;
sin_rom[896] = 2121;
sin_rom[897] = 2095;
sin_rom[898] = 2070;
sin_rom[899] = 2044;
sin_rom[900] = 2019;
sin_rom[901] = 1993;
sin_rom[902] = 1968;
sin_rom[903] = 1942;
sin_rom[904] = 1917;
sin_rom[905] = 1891;
sin_rom[906] = 1865;
sin_rom[907] = 1840;
sin_rom[908] = 1814;
sin_rom[909] = 1788;
sin_rom[910] = 1763;
sin_rom[911] = 1737;
sin_rom[912] = 1711;
sin_rom[913] = 1685;
sin_rom[914] = 1660;
sin_rom[915] = 1634;
sin_rom[916] = 1608;
sin_rom[917] = 1582;
sin_rom[918] = 1556;
sin_rom[919] = 1531;
sin_rom[920] = 1505;
sin_rom[921] = 1479;
sin_rom[922] = 1453;
sin_rom[923] = 1427;
sin_rom[924] = 1401;
sin_rom[925] = 1375;
sin_rom[926] = 1349;
sin_rom[927] = 1323;
sin_rom[928] = 1297;
sin_rom[929] = 1271;
sin_rom[930] = 1245;
sin_rom[931] = 1219;
sin_rom[932] = 1193;
sin_rom[933] = 1167;
sin_rom[934] = 1141;
sin_rom[935] = 1115;
sin_rom[936] = 1089;
sin_rom[937] = 1063;
sin_rom[938] = 1037;
sin_rom[939] = 1010;
sin_rom[940] = 984;
sin_rom[941] = 958;
sin_rom[942] = 932;
sin_rom[943] = 906;
sin_rom[944] = 880;
sin_rom[945] = 854;
sin_rom[946] = 827;
sin_rom[947] = 801;
sin_rom[948] = 775;
sin_rom[949] = 749;
sin_rom[950] = 722;
sin_rom[951] = 696;
sin_rom[952] = 670;
sin_rom[953] = 644;
sin_rom[954] = 618;
sin_rom[955] = 591;
sin_rom[956] = 565;
sin_rom[957] = 539;
sin_rom[958] = 512;
sin_rom[959] = 486;
sin_rom[960] = 460;
sin_rom[961] = 434;
sin_rom[962] = 407;
sin_rom[963] = 381;
sin_rom[964] = 355;
sin_rom[965] = 328;
sin_rom[966] = 302;
sin_rom[967] = 276;
sin_rom[968] = 249;
sin_rom[969] = 223;
sin_rom[970] = 197;
sin_rom[971] = 171;
sin_rom[972] = 144;
sin_rom[973] = 118;
sin_rom[974] = 92;
sin_rom[975] = 65;
sin_rom[976] = 39;
sin_rom[977] = 13;
sin_rom[978] = -13;
sin_rom[979] = -39;
sin_rom[980] = -65;
sin_rom[981] = -92;
sin_rom[982] = -118;
sin_rom[983] = -144;
sin_rom[984] = -171;
sin_rom[985] = -197;
sin_rom[986] = -223;
sin_rom[987] = -250;
sin_rom[988] = -276;
sin_rom[989] = -302;
sin_rom[990] = -329;
sin_rom[991] = -355;
sin_rom[992] = -381;
sin_rom[993] = -408;
sin_rom[994] = -434;
sin_rom[995] = -460;
sin_rom[996] = -486;
sin_rom[997] = -513;
sin_rom[998] = -539;
sin_rom[999] = -565;
sin_rom[1000] = -591;
sin_rom[1001] = -618;
sin_rom[1002] = -644;
sin_rom[1003] = -670;
sin_rom[1004] = -696;
sin_rom[1005] = -723;
sin_rom[1006] = -749;
sin_rom[1007] = -775;
sin_rom[1008] = -801;
sin_rom[1009] = -828;
sin_rom[1010] = -854;
sin_rom[1011] = -880;
sin_rom[1012] = -906;
sin_rom[1013] = -932;
sin_rom[1014] = -958;
sin_rom[1015] = -985;
sin_rom[1016] = -1011;
sin_rom[1017] = -1037;
sin_rom[1018] = -1063;
sin_rom[1019] = -1089;
sin_rom[1020] = -1115;
sin_rom[1021] = -1141;
sin_rom[1022] = -1167;
sin_rom[1023] = -1193;
sin_rom[1024] = -1219;
sin_rom[1025] = -1245;
sin_rom[1026] = -1271;
sin_rom[1027] = -1297;
sin_rom[1028] = -1323;
sin_rom[1029] = -1349;
sin_rom[1030] = -1375;
sin_rom[1031] = -1401;
sin_rom[1032] = -1427;
sin_rom[1033] = -1453;
sin_rom[1034] = -1479;
sin_rom[1035] = -1505;
sin_rom[1036] = -1531;
sin_rom[1037] = -1557;
sin_rom[1038] = -1582;
sin_rom[1039] = -1608;
sin_rom[1040] = -1634;
sin_rom[1041] = -1660;
sin_rom[1042] = -1686;
sin_rom[1043] = -1711;
sin_rom[1044] = -1737;
sin_rom[1045] = -1763;
sin_rom[1046] = -1789;
sin_rom[1047] = -1814;
sin_rom[1048] = -1840;
sin_rom[1049] = -1866;
sin_rom[1050] = -1891;
sin_rom[1051] = -1917;
sin_rom[1052] = -1942;
sin_rom[1053] = -1968;
sin_rom[1054] = -1994;
sin_rom[1055] = -2019;
sin_rom[1056] = -2045;
sin_rom[1057] = -2070;
sin_rom[1058] = -2095;
sin_rom[1059] = -2121;
sin_rom[1060] = -2146;
sin_rom[1061] = -2172;
sin_rom[1062] = -2197;
sin_rom[1063] = -2222;
sin_rom[1064] = -2248;
sin_rom[1065] = -2273;
sin_rom[1066] = -2298;
sin_rom[1067] = -2324;
sin_rom[1068] = -2349;
sin_rom[1069] = -2374;
sin_rom[1070] = -2399;
sin_rom[1071] = -2424;
sin_rom[1072] = -2450;
sin_rom[1073] = -2475;
sin_rom[1074] = -2500;
sin_rom[1075] = -2525;
sin_rom[1076] = -2550;
sin_rom[1077] = -2575;
sin_rom[1078] = -2600;
sin_rom[1079] = -2625;
sin_rom[1080] = -2650;
sin_rom[1081] = -2675;
sin_rom[1082] = -2699;
sin_rom[1083] = -2724;
sin_rom[1084] = -2749;
sin_rom[1085] = -2774;
sin_rom[1086] = -2799;
sin_rom[1087] = -2823;
sin_rom[1088] = -2848;
sin_rom[1089] = -2873;
sin_rom[1090] = -2897;
sin_rom[1091] = -2922;
sin_rom[1092] = -2947;
sin_rom[1093] = -2971;
sin_rom[1094] = -2996;
sin_rom[1095] = -3020;
sin_rom[1096] = -3045;
sin_rom[1097] = -3069;
sin_rom[1098] = -3093;
sin_rom[1099] = -3118;
sin_rom[1100] = -3142;
sin_rom[1101] = -3166;
sin_rom[1102] = -3191;
sin_rom[1103] = -3215;
sin_rom[1104] = -3239;
sin_rom[1105] = -3263;
sin_rom[1106] = -3287;
sin_rom[1107] = -3312;
sin_rom[1108] = -3336;
sin_rom[1109] = -3360;
sin_rom[1110] = -3384;
sin_rom[1111] = -3408;
sin_rom[1112] = -3432;
sin_rom[1113] = -3455;
sin_rom[1114] = -3479;
sin_rom[1115] = -3503;
sin_rom[1116] = -3527;
sin_rom[1117] = -3551;
sin_rom[1118] = -3574;
sin_rom[1119] = -3598;
sin_rom[1120] = -3622;
sin_rom[1121] = -3645;
sin_rom[1122] = -3669;
sin_rom[1123] = -3692;
sin_rom[1124] = -3716;
sin_rom[1125] = -3739;
sin_rom[1126] = -3763;
sin_rom[1127] = -3786;
sin_rom[1128] = -3809;
sin_rom[1129] = -3833;
sin_rom[1130] = -3856;
sin_rom[1131] = -3879;
sin_rom[1132] = -3902;
sin_rom[1133] = -3925;
sin_rom[1134] = -3948;
sin_rom[1135] = -3971;
sin_rom[1136] = -3995;
sin_rom[1137] = -4017;
sin_rom[1138] = -4040;
sin_rom[1139] = -4063;
sin_rom[1140] = -4086;
sin_rom[1141] = -4109;
sin_rom[1142] = -4132;
sin_rom[1143] = -4154;
sin_rom[1144] = -4177;
sin_rom[1145] = -4200;
sin_rom[1146] = -4222;
sin_rom[1147] = -4245;
sin_rom[1148] = -4267;
sin_rom[1149] = -4290;
sin_rom[1150] = -4312;
sin_rom[1151] = -4335;
sin_rom[1152] = -4357;
sin_rom[1153] = -4379;
sin_rom[1154] = -4401;
sin_rom[1155] = -4424;
sin_rom[1156] = -4446;
sin_rom[1157] = -4468;
sin_rom[1158] = -4490;
sin_rom[1159] = -4512;
sin_rom[1160] = -4534;
sin_rom[1161] = -4556;
sin_rom[1162] = -4577;
sin_rom[1163] = -4599;
sin_rom[1164] = -4621;
sin_rom[1165] = -4643;
sin_rom[1166] = -4664;
sin_rom[1167] = -4686;
sin_rom[1168] = -4708;
sin_rom[1169] = -4729;
sin_rom[1170] = -4751;
sin_rom[1171] = -4772;
sin_rom[1172] = -4793;
sin_rom[1173] = -4815;
sin_rom[1174] = -4836;
sin_rom[1175] = -4857;
sin_rom[1176] = -4878;
sin_rom[1177] = -4900;
sin_rom[1178] = -4921;
sin_rom[1179] = -4942;
sin_rom[1180] = -4963;
sin_rom[1181] = -4984;
sin_rom[1182] = -5004;
sin_rom[1183] = -5025;
sin_rom[1184] = -5046;
sin_rom[1185] = -5067;
sin_rom[1186] = -5087;
sin_rom[1187] = -5108;
sin_rom[1188] = -5129;
sin_rom[1189] = -5149;
sin_rom[1190] = -5169;
sin_rom[1191] = -5190;
sin_rom[1192] = -5210;
sin_rom[1193] = -5231;
sin_rom[1194] = -5251;
sin_rom[1195] = -5271;
sin_rom[1196] = -5291;
sin_rom[1197] = -5311;
sin_rom[1198] = -5331;
sin_rom[1199] = -5351;
sin_rom[1200] = -5371;
sin_rom[1201] = -5391;
sin_rom[1202] = -5411;
sin_rom[1203] = -5430;
sin_rom[1204] = -5450;
sin_rom[1205] = -5470;
sin_rom[1206] = -5489;
sin_rom[1207] = -5509;
sin_rom[1208] = -5528;
sin_rom[1209] = -5548;
sin_rom[1210] = -5567;
sin_rom[1211] = -5586;
sin_rom[1212] = -5605;
sin_rom[1213] = -5625;
sin_rom[1214] = -5644;
sin_rom[1215] = -5663;
sin_rom[1216] = -5682;
sin_rom[1217] = -5701;
sin_rom[1218] = -5720;
sin_rom[1219] = -5738;
sin_rom[1220] = -5757;
sin_rom[1221] = -5776;
sin_rom[1222] = -5795;
sin_rom[1223] = -5813;
sin_rom[1224] = -5832;
sin_rom[1225] = -5850;
sin_rom[1226] = -5869;
sin_rom[1227] = -5887;
sin_rom[1228] = -5905;
sin_rom[1229] = -5923;
sin_rom[1230] = -5941;
sin_rom[1231] = -5960;
sin_rom[1232] = -5978;
sin_rom[1233] = -5996;
sin_rom[1234] = -6013;
sin_rom[1235] = -6031;
sin_rom[1236] = -6049;
sin_rom[1237] = -6067;
sin_rom[1238] = -6085;
sin_rom[1239] = -6102;
sin_rom[1240] = -6120;
sin_rom[1241] = -6137;
sin_rom[1242] = -6155;
sin_rom[1243] = -6172;
sin_rom[1244] = -6189;
sin_rom[1245] = -6206;
sin_rom[1246] = -6223;
sin_rom[1247] = -6241;
sin_rom[1248] = -6258;
sin_rom[1249] = -6275;
sin_rom[1250] = -6291;
sin_rom[1251] = -6308;
sin_rom[1252] = -6325;
sin_rom[1253] = -6342;
sin_rom[1254] = -6358;
sin_rom[1255] = -6375;
sin_rom[1256] = -6391;
sin_rom[1257] = -6408;
sin_rom[1258] = -6424;
sin_rom[1259] = -6441;
sin_rom[1260] = -6457;
sin_rom[1261] = -6473;
sin_rom[1262] = -6489;
sin_rom[1263] = -6505;
sin_rom[1264] = -6521;
sin_rom[1265] = -6537;
sin_rom[1266] = -6553;
sin_rom[1267] = -6569;
sin_rom[1268] = -6584;
sin_rom[1269] = -6600;
sin_rom[1270] = -6615;
sin_rom[1271] = -6631;
sin_rom[1272] = -6646;
sin_rom[1273] = -6662;
sin_rom[1274] = -6677;
sin_rom[1275] = -6692;
sin_rom[1276] = -6707;
sin_rom[1277] = -6722;
sin_rom[1278] = -6737;
sin_rom[1279] = -6752;
sin_rom[1280] = -6767;
sin_rom[1281] = -6782;
sin_rom[1282] = -6797;
sin_rom[1283] = -6811;
sin_rom[1284] = -6826;
sin_rom[1285] = -6841;
sin_rom[1286] = -6855;
sin_rom[1287] = -6869;
sin_rom[1288] = -6884;
sin_rom[1289] = -6898;
sin_rom[1290] = -6912;
sin_rom[1291] = -6926;
sin_rom[1292] = -6940;
sin_rom[1293] = -6954;
sin_rom[1294] = -6968;
sin_rom[1295] = -6982;
sin_rom[1296] = -6996;
sin_rom[1297] = -7009;
sin_rom[1298] = -7023;
sin_rom[1299] = -7036;
sin_rom[1300] = -7050;
sin_rom[1301] = -7063;
sin_rom[1302] = -7076;
sin_rom[1303] = -7090;
sin_rom[1304] = -7103;
sin_rom[1305] = -7116;
sin_rom[1306] = -7129;
sin_rom[1307] = -7142;
sin_rom[1308] = -7155;
sin_rom[1309] = -7167;
sin_rom[1310] = -7180;
sin_rom[1311] = -7193;
sin_rom[1312] = -7205;
sin_rom[1313] = -7218;
sin_rom[1314] = -7230;
sin_rom[1315] = -7243;
sin_rom[1316] = -7255;
sin_rom[1317] = -7267;
sin_rom[1318] = -7279;
sin_rom[1319] = -7291;
sin_rom[1320] = -7303;
sin_rom[1321] = -7315;
sin_rom[1322] = -7327;
sin_rom[1323] = -7339;
sin_rom[1324] = -7350;
sin_rom[1325] = -7362;
sin_rom[1326] = -7373;
sin_rom[1327] = -7385;
sin_rom[1328] = -7396;
sin_rom[1329] = -7407;
sin_rom[1330] = -7419;
sin_rom[1331] = -7430;
sin_rom[1332] = -7441;
sin_rom[1333] = -7452;
sin_rom[1334] = -7463;
sin_rom[1335] = -7473;
sin_rom[1336] = -7484;
sin_rom[1337] = -7495;
sin_rom[1338] = -7505;
sin_rom[1339] = -7516;
sin_rom[1340] = -7526;
sin_rom[1341] = -7537;
sin_rom[1342] = -7547;
sin_rom[1343] = -7557;
sin_rom[1344] = -7567;
sin_rom[1345] = -7577;
sin_rom[1346] = -7587;
sin_rom[1347] = -7597;
sin_rom[1348] = -7607;
sin_rom[1349] = -7617;
sin_rom[1350] = -7626;
sin_rom[1351] = -7636;
sin_rom[1352] = -7645;
sin_rom[1353] = -7655;
sin_rom[1354] = -7664;
sin_rom[1355] = -7673;
sin_rom[1356] = -7683;
sin_rom[1357] = -7692;
sin_rom[1358] = -7701;
sin_rom[1359] = -7710;
sin_rom[1360] = -7719;
sin_rom[1361] = -7727;
sin_rom[1362] = -7736;
sin_rom[1363] = -7745;
sin_rom[1364] = -7753;
sin_rom[1365] = -7762;
sin_rom[1366] = -7770;
sin_rom[1367] = -7778;
sin_rom[1368] = -7787;
sin_rom[1369] = -7795;
sin_rom[1370] = -7803;
sin_rom[1371] = -7811;
sin_rom[1372] = -7819;
sin_rom[1373] = -7826;
sin_rom[1374] = -7834;
sin_rom[1375] = -7842;
sin_rom[1376] = -7849;
sin_rom[1377] = -7857;
sin_rom[1378] = -7864;
sin_rom[1379] = -7872;
sin_rom[1380] = -7879;
sin_rom[1381] = -7886;
sin_rom[1382] = -7893;
sin_rom[1383] = -7900;
sin_rom[1384] = -7907;
sin_rom[1385] = -7914;
sin_rom[1386] = -7921;
sin_rom[1387] = -7927;
sin_rom[1388] = -7934;
sin_rom[1389] = -7940;
sin_rom[1390] = -7947;
sin_rom[1391] = -7953;
sin_rom[1392] = -7959;
sin_rom[1393] = -7966;
sin_rom[1394] = -7972;
sin_rom[1395] = -7978;
sin_rom[1396] = -7984;
sin_rom[1397] = -7989;
sin_rom[1398] = -7995;
sin_rom[1399] = -8001;
sin_rom[1400] = -8007;
sin_rom[1401] = -8012;
sin_rom[1402] = -8018;
sin_rom[1403] = -8023;
sin_rom[1404] = -8028;
sin_rom[1405] = -8033;
sin_rom[1406] = -8038;
sin_rom[1407] = -8043;
sin_rom[1408] = -8048;
sin_rom[1409] = -8053;
sin_rom[1410] = -8058;
sin_rom[1411] = -8063;
sin_rom[1412] = -8067;
sin_rom[1413] = -8072;
sin_rom[1414] = -8076;
sin_rom[1415] = -8081;
sin_rom[1416] = -8085;
sin_rom[1417] = -8089;
sin_rom[1418] = -8093;
sin_rom[1419] = -8097;
sin_rom[1420] = -8101;
sin_rom[1421] = -8105;
sin_rom[1422] = -8109;
sin_rom[1423] = -8113;
sin_rom[1424] = -8116;
sin_rom[1425] = -8120;
sin_rom[1426] = -8123;
sin_rom[1427] = -8126;
sin_rom[1428] = -8130;
sin_rom[1429] = -8133;
sin_rom[1430] = -8136;
sin_rom[1431] = -8139;
sin_rom[1432] = -8142;
sin_rom[1433] = -8145;
sin_rom[1434] = -8148;
sin_rom[1435] = -8150;
sin_rom[1436] = -8153;
sin_rom[1437] = -8155;
sin_rom[1438] = -8158;
sin_rom[1439] = -8160;
sin_rom[1440] = -8162;
sin_rom[1441] = -8165;
sin_rom[1442] = -8167;
sin_rom[1443] = -8169;
sin_rom[1444] = -8171;
sin_rom[1445] = -8172;
sin_rom[1446] = -8174;
sin_rom[1447] = -8176;
sin_rom[1448] = -8177;
sin_rom[1449] = -8179;
sin_rom[1450] = -8180;
sin_rom[1451] = -8182;
sin_rom[1452] = -8183;
sin_rom[1453] = -8184;
sin_rom[1454] = -8185;
sin_rom[1455] = -8186;
sin_rom[1456] = -8187;
sin_rom[1457] = -8188;
sin_rom[1458] = -8189;
sin_rom[1459] = -8189;
sin_rom[1460] = -8190;
sin_rom[1461] = -8190;
sin_rom[1462] = -8191;
sin_rom[1463] = -8191;
sin_rom[1464] = -8191;
sin_rom[1465] = -8191;
sin_rom[1466] = -8191;
sin_rom[1467] = -8191;
sin_rom[1468] = -8191;
sin_rom[1469] = -8191;
sin_rom[1470] = -8191;
sin_rom[1471] = -8191;
sin_rom[1472] = -8190;
sin_rom[1473] = -8190;
sin_rom[1474] = -8189;
sin_rom[1475] = -8188;
sin_rom[1476] = -8187;
sin_rom[1477] = -8187;
sin_rom[1478] = -8186;
sin_rom[1479] = -8185;
sin_rom[1480] = -8183;
sin_rom[1481] = -8182;
sin_rom[1482] = -8181;
sin_rom[1483] = -8180;
sin_rom[1484] = -8178;
sin_rom[1485] = -8177;
sin_rom[1486] = -8175;
sin_rom[1487] = -8173;
sin_rom[1488] = -8171;
sin_rom[1489] = -8170;
sin_rom[1490] = -8168;
sin_rom[1491] = -8166;
sin_rom[1492] = -8163;
sin_rom[1493] = -8161;
sin_rom[1494] = -8159;
sin_rom[1495] = -8157;
sin_rom[1496] = -8154;
sin_rom[1497] = -8152;
sin_rom[1498] = -8149;
sin_rom[1499] = -8146;
sin_rom[1500] = -8143;
sin_rom[1501] = -8140;
sin_rom[1502] = -8137;
sin_rom[1503] = -8134;
sin_rom[1504] = -8131;
sin_rom[1505] = -8128;
sin_rom[1506] = -8125;
sin_rom[1507] = -8121;
sin_rom[1508] = -8118;
sin_rom[1509] = -8114;
sin_rom[1510] = -8111;
sin_rom[1511] = -8107;
sin_rom[1512] = -8103;
sin_rom[1513] = -8099;
sin_rom[1514] = -8095;
sin_rom[1515] = -8091;
sin_rom[1516] = -8087;
sin_rom[1517] = -8083;
sin_rom[1518] = -8078;
sin_rom[1519] = -8074;
sin_rom[1520] = -8070;
sin_rom[1521] = -8065;
sin_rom[1522] = -8060;
sin_rom[1523] = -8056;
sin_rom[1524] = -8051;
sin_rom[1525] = -8046;
sin_rom[1526] = -8041;
sin_rom[1527] = -8036;
sin_rom[1528] = -8031;
sin_rom[1529] = -8025;
sin_rom[1530] = -8020;
sin_rom[1531] = -8015;
sin_rom[1532] = -8009;
sin_rom[1533] = -8004;
sin_rom[1534] = -7998;
sin_rom[1535] = -7992;
sin_rom[1536] = -7986;
sin_rom[1537] = -7981;
sin_rom[1538] = -7975;
sin_rom[1539] = -7969;
sin_rom[1540] = -7962;
sin_rom[1541] = -7956;
sin_rom[1542] = -7950;
sin_rom[1543] = -7943;
sin_rom[1544] = -7937;
sin_rom[1545] = -7930;
sin_rom[1546] = -7924;
sin_rom[1547] = -7917;
sin_rom[1548] = -7910;
sin_rom[1549] = -7903;
sin_rom[1550] = -7896;
sin_rom[1551] = -7889;
sin_rom[1552] = -7882;
sin_rom[1553] = -7875;
sin_rom[1554] = -7868;
sin_rom[1555] = -7860;
sin_rom[1556] = -7853;
sin_rom[1557] = -7845;
sin_rom[1558] = -7838;
sin_rom[1559] = -7830;
sin_rom[1560] = -7822;
sin_rom[1561] = -7815;
sin_rom[1562] = -7807;
sin_rom[1563] = -7799;
sin_rom[1564] = -7790;
sin_rom[1565] = -7782;
sin_rom[1566] = -7774;
sin_rom[1567] = -7766;
sin_rom[1568] = -7757;
sin_rom[1569] = -7749;
sin_rom[1570] = -7740;
sin_rom[1571] = -7732;
sin_rom[1572] = -7723;
sin_rom[1573] = -7714;
sin_rom[1574] = -7705;
sin_rom[1575] = -7696;
sin_rom[1576] = -7687;
sin_rom[1577] = -7678;
sin_rom[1578] = -7669;
sin_rom[1579] = -7659;
sin_rom[1580] = -7650;
sin_rom[1581] = -7641;
sin_rom[1582] = -7631;
sin_rom[1583] = -7621;
sin_rom[1584] = -7612;
sin_rom[1585] = -7602;
sin_rom[1586] = -7592;
sin_rom[1587] = -7582;
sin_rom[1588] = -7572;
sin_rom[1589] = -7562;
sin_rom[1590] = -7552;
sin_rom[1591] = -7542;
sin_rom[1592] = -7531;
sin_rom[1593] = -7521;
sin_rom[1594] = -7511;
sin_rom[1595] = -7500;
sin_rom[1596] = -7489;
sin_rom[1597] = -7479;
sin_rom[1598] = -7468;
sin_rom[1599] = -7457;
sin_rom[1600] = -7446;
sin_rom[1601] = -7435;
sin_rom[1602] = -7424;
sin_rom[1603] = -7413;
sin_rom[1604] = -7402;
sin_rom[1605] = -7390;
sin_rom[1606] = -7379;
sin_rom[1607] = -7367;
sin_rom[1608] = -7356;
sin_rom[1609] = -7344;
sin_rom[1610] = -7333;
sin_rom[1611] = -7321;
sin_rom[1612] = -7309;
sin_rom[1613] = -7297;
sin_rom[1614] = -7285;
sin_rom[1615] = -7273;
sin_rom[1616] = -7261;
sin_rom[1617] = -7249;
sin_rom[1618] = -7236;
sin_rom[1619] = -7224;
sin_rom[1620] = -7211;
sin_rom[1621] = -7199;
sin_rom[1622] = -7186;
sin_rom[1623] = -7174;
sin_rom[1624] = -7161;
sin_rom[1625] = -7148;
sin_rom[1626] = -7135;
sin_rom[1627] = -7122;
sin_rom[1628] = -7109;
sin_rom[1629] = -7096;
sin_rom[1630] = -7083;
sin_rom[1631] = -7070;
sin_rom[1632] = -7056;
sin_rom[1633] = -7043;
sin_rom[1634] = -7029;
sin_rom[1635] = -7016;
sin_rom[1636] = -7002;
sin_rom[1637] = -6989;
sin_rom[1638] = -6975;
sin_rom[1639] = -6961;
sin_rom[1640] = -6947;
sin_rom[1641] = -6933;
sin_rom[1642] = -6919;
sin_rom[1643] = -6905;
sin_rom[1644] = -6891;
sin_rom[1645] = -6876;
sin_rom[1646] = -6862;
sin_rom[1647] = -6848;
sin_rom[1648] = -6833;
sin_rom[1649] = -6819;
sin_rom[1650] = -6804;
sin_rom[1651] = -6789;
sin_rom[1652] = -6774;
sin_rom[1653] = -6760;
sin_rom[1654] = -6745;
sin_rom[1655] = -6730;
sin_rom[1656] = -6715;
sin_rom[1657] = -6700;
sin_rom[1658] = -6684;
sin_rom[1659] = -6669;
sin_rom[1660] = -6654;
sin_rom[1661] = -6638;
sin_rom[1662] = -6623;
sin_rom[1663] = -6607;
sin_rom[1664] = -6592;
sin_rom[1665] = -6576;
sin_rom[1666] = -6560;
sin_rom[1667] = -6545;
sin_rom[1668] = -6529;
sin_rom[1669] = -6513;
sin_rom[1670] = -6497;
sin_rom[1671] = -6481;
sin_rom[1672] = -6465;
sin_rom[1673] = -6448;
sin_rom[1674] = -6432;
sin_rom[1675] = -6416;
sin_rom[1676] = -6399;
sin_rom[1677] = -6383;
sin_rom[1678] = -6366;
sin_rom[1679] = -6350;
sin_rom[1680] = -6333;
sin_rom[1681] = -6316;
sin_rom[1682] = -6300;
sin_rom[1683] = -6283;
sin_rom[1684] = -6266;
sin_rom[1685] = -6249;
sin_rom[1686] = -6232;
sin_rom[1687] = -6215;
sin_rom[1688] = -6198;
sin_rom[1689] = -6180;
sin_rom[1690] = -6163;
sin_rom[1691] = -6146;
sin_rom[1692] = -6128;
sin_rom[1693] = -6111;
sin_rom[1694] = -6093;
sin_rom[1695] = -6075;
sin_rom[1696] = -6058;
sin_rom[1697] = -6040;
sin_rom[1698] = -6022;
sin_rom[1699] = -6004;
sin_rom[1700] = -5986;
sin_rom[1701] = -5968;
sin_rom[1702] = -5950;
sin_rom[1703] = -5932;
sin_rom[1704] = -5914;
sin_rom[1705] = -5896;
sin_rom[1706] = -5877;
sin_rom[1707] = -5859;
sin_rom[1708] = -5841;
sin_rom[1709] = -5822;
sin_rom[1710] = -5804;
sin_rom[1711] = -5785;
sin_rom[1712] = -5766;
sin_rom[1713] = -5748;
sin_rom[1714] = -5729;
sin_rom[1715] = -5710;
sin_rom[1716] = -5691;
sin_rom[1717] = -5672;
sin_rom[1718] = -5653;
sin_rom[1719] = -5634;
sin_rom[1720] = -5615;
sin_rom[1721] = -5596;
sin_rom[1722] = -5576;
sin_rom[1723] = -5557;
sin_rom[1724] = -5538;
sin_rom[1725] = -5518;
sin_rom[1726] = -5499;
sin_rom[1727] = -5479;
sin_rom[1728] = -5460;
sin_rom[1729] = -5440;
sin_rom[1730] = -5420;
sin_rom[1731] = -5400;
sin_rom[1732] = -5381;
sin_rom[1733] = -5361;
sin_rom[1734] = -5341;
sin_rom[1735] = -5321;
sin_rom[1736] = -5301;
sin_rom[1737] = -5281;
sin_rom[1738] = -5261;
sin_rom[1739] = -5240;
sin_rom[1740] = -5220;
sin_rom[1741] = -5200;
sin_rom[1742] = -5179;
sin_rom[1743] = -5159;
sin_rom[1744] = -5139;
sin_rom[1745] = -5118;
sin_rom[1746] = -5097;
sin_rom[1747] = -5077;
sin_rom[1748] = -5056;
sin_rom[1749] = -5035;
sin_rom[1750] = -5015;
sin_rom[1751] = -4994;
sin_rom[1752] = -4973;
sin_rom[1753] = -4952;
sin_rom[1754] = -4931;
sin_rom[1755] = -4910;
sin_rom[1756] = -4889;
sin_rom[1757] = -4868;
sin_rom[1758] = -4846;
sin_rom[1759] = -4825;
sin_rom[1760] = -4804;
sin_rom[1761] = -4782;
sin_rom[1762] = -4761;
sin_rom[1763] = -4740;
sin_rom[1764] = -4718;
sin_rom[1765] = -4697;
sin_rom[1766] = -4675;
sin_rom[1767] = -4653;
sin_rom[1768] = -4632;
sin_rom[1769] = -4610;
sin_rom[1770] = -4588;
sin_rom[1771] = -4566;
sin_rom[1772] = -4544;
sin_rom[1773] = -4522;
sin_rom[1774] = -4500;
sin_rom[1775] = -4478;
sin_rom[1776] = -4456;
sin_rom[1777] = -4434;
sin_rom[1778] = -4412;
sin_rom[1779] = -4390;
sin_rom[1780] = -4368;
sin_rom[1781] = -4345;
sin_rom[1782] = -4323;
sin_rom[1783] = -4301;
sin_rom[1784] = -4278;
sin_rom[1785] = -4256;
sin_rom[1786] = -4233;
sin_rom[1787] = -4211;
sin_rom[1788] = -4188;
sin_rom[1789] = -4165;
sin_rom[1790] = -4143;
sin_rom[1791] = -4120;
sin_rom[1792] = -4097;
sin_rom[1793] = -4074;
sin_rom[1794] = -4052;
sin_rom[1795] = -4029;
sin_rom[1796] = -4006;
sin_rom[1797] = -3983;
sin_rom[1798] = -3960;
sin_rom[1799] = -3937;
sin_rom[1800] = -3913;
sin_rom[1801] = -3890;
sin_rom[1802] = -3867;
sin_rom[1803] = -3844;
sin_rom[1804] = -3821;
sin_rom[1805] = -3797;
sin_rom[1806] = -3774;
sin_rom[1807] = -3751;
sin_rom[1808] = -3727;
sin_rom[1809] = -3704;
sin_rom[1810] = -3680;
sin_rom[1811] = -3657;
sin_rom[1812] = -3633;
sin_rom[1813] = -3609;
sin_rom[1814] = -3586;
sin_rom[1815] = -3562;
sin_rom[1816] = -3538;
sin_rom[1817] = -3515;
sin_rom[1818] = -3491;
sin_rom[1819] = -3467;
sin_rom[1820] = -3443;
sin_rom[1821] = -3419;
sin_rom[1822] = -3395;
sin_rom[1823] = -3371;
sin_rom[1824] = -3347;
sin_rom[1825] = -3323;
sin_rom[1826] = -3299;
sin_rom[1827] = -3275;
sin_rom[1828] = -3251;
sin_rom[1829] = -3227;
sin_rom[1830] = -3203;
sin_rom[1831] = -3178;
sin_rom[1832] = -3154;
sin_rom[1833] = -3130;
sin_rom[1834] = -3105;
sin_rom[1835] = -3081;
sin_rom[1836] = -3057;
sin_rom[1837] = -3032;
sin_rom[1838] = -3008;
sin_rom[1839] = -2983;
sin_rom[1840] = -2959;
sin_rom[1841] = -2934;
sin_rom[1842] = -2909;
sin_rom[1843] = -2885;
sin_rom[1844] = -2860;
sin_rom[1845] = -2835;
sin_rom[1846] = -2811;
sin_rom[1847] = -2786;
sin_rom[1848] = -2761;
sin_rom[1849] = -2736;
sin_rom[1850] = -2712;
sin_rom[1851] = -2687;
sin_rom[1852] = -2662;
sin_rom[1853] = -2637;
sin_rom[1854] = -2612;
sin_rom[1855] = -2587;
sin_rom[1856] = -2562;
sin_rom[1857] = -2537;
sin_rom[1858] = -2512;
sin_rom[1859] = -2487;
sin_rom[1860] = -2462;
sin_rom[1861] = -2437;
sin_rom[1862] = -2412;
sin_rom[1863] = -2386;
sin_rom[1864] = -2361;
sin_rom[1865] = -2336;
sin_rom[1866] = -2311;
sin_rom[1867] = -2285;
sin_rom[1868] = -2260;
sin_rom[1869] = -2235;
sin_rom[1870] = -2209;
sin_rom[1871] = -2184;
sin_rom[1872] = -2159;
sin_rom[1873] = -2133;
sin_rom[1874] = -2108;
sin_rom[1875] = -2082;
sin_rom[1876] = -2057;
sin_rom[1877] = -2031;
sin_rom[1878] = -2006;
sin_rom[1879] = -1980;
sin_rom[1880] = -1955;
sin_rom[1881] = -1929;
sin_rom[1882] = -1904;
sin_rom[1883] = -1878;
sin_rom[1884] = -1852;
sin_rom[1885] = -1827;
sin_rom[1886] = -1801;
sin_rom[1887] = -1775;
sin_rom[1888] = -1750;
sin_rom[1889] = -1724;
sin_rom[1890] = -1698;
sin_rom[1891] = -1672;
sin_rom[1892] = -1647;
sin_rom[1893] = -1621;
sin_rom[1894] = -1595;
sin_rom[1895] = -1569;
sin_rom[1896] = -1543;
sin_rom[1897] = -1517;
sin_rom[1898] = -1492;
sin_rom[1899] = -1466;
sin_rom[1900] = -1440;
sin_rom[1901] = -1414;
sin_rom[1902] = -1388;
sin_rom[1903] = -1362;
sin_rom[1904] = -1336;
sin_rom[1905] = -1310;
sin_rom[1906] = -1284;
sin_rom[1907] = -1258;
sin_rom[1908] = -1232;
sin_rom[1909] = -1206;
sin_rom[1910] = -1180;
sin_rom[1911] = -1154;
sin_rom[1912] = -1128;
sin_rom[1913] = -1102;
sin_rom[1914] = -1076;
sin_rom[1915] = -1050;
sin_rom[1916] = -1023;
sin_rom[1917] = -997;
sin_rom[1918] = -971;
sin_rom[1919] = -945;
sin_rom[1920] = -919;
sin_rom[1921] = -893;
sin_rom[1922] = -866;
sin_rom[1923] = -840;
sin_rom[1924] = -814;
sin_rom[1925] = -788;
sin_rom[1926] = -762;
sin_rom[1927] = -735;
sin_rom[1928] = -709;
sin_rom[1929] = -683;
sin_rom[1930] = -657;
sin_rom[1931] = -631;
sin_rom[1932] = -604;
sin_rom[1933] = -578;
sin_rom[1934] = -552;
sin_rom[1935] = -525;
sin_rom[1936] = -499;
sin_rom[1937] = -473;
sin_rom[1938] = -447;
sin_rom[1939] = -420;
sin_rom[1940] = -394;
sin_rom[1941] = -368;
sin_rom[1942] = -341;
sin_rom[1943] = -315;
sin_rom[1944] = -289;
sin_rom[1945] = -263;
sin_rom[1946] = -236;
sin_rom[1947] = -210;
sin_rom[1948] = -184;
sin_rom[1949] = -157;
sin_rom[1950] = -131;
sin_rom[1951] = -105;
sin_rom[1952] = -78;
sin_rom[1953] = -52;
end


reg [18:0]addr = 0;
reg [18:0]addr_r;

always@(posedge clk)begin
    if(addr+freq<500000)
        addr<=addr+freq;
    else
        addr<=addr+freq-500000;
    if(addr+phase<500000)
        addr_r<=addr+phase;
    else
        addr<=addr+phase-500000;
    dds_o<=sin_rom[addr_r[18:8]];
end

endmodule